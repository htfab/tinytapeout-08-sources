** sch_path: /home/ttuser/test0/tt08-bgr/xschem/opamp_l_pl.sch
**.subckt opamp_l_pl
x1 VDD VSS in MINUS PLUS out opamp_l
V1 VDD GND 1.8
V2 VSS GND 0
I0 VDD in 37.545u
V5 MINUS GND 0.75
V6 PLUS MINUS dc 0 ac 1 0
.save v(out)
x2 VDD VSS in MINUS PLUS outr opamp_l_parax
.save v(outr)
C1 out GND 1p m=1
C2 outr GND 1p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




.option savecurrents
.control
  save all
  ac dec 20 1k 2G
  remzerovec
  write opamp_l.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  opamp_l.sym # of pins=6
** sym_path: /home/ttuser/test0/tt08-bgr/xschem/opamp_l.sym
** sch_path: /home/ttuser/test0/tt08-bgr/xschem/opamp_l.sch
.subckt opamp_l VDD VSS in MINUS PLUS opout
*.ipin VDD
*.ipin VSS
*.ipin in
*.ipin MINUS
*.ipin PLUS
*.iopin opout
XM4 opout MINUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 PLUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 opout net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net1 in VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 in in VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  opamp_l_parax.sym # of pins=6
** sym_path: /home/ttuser/test0/tt08-bgr/xschem/opamp_l.sym
.include /home/ttuser/test0/tt08-bgr/mag/opamp_l.sim.spice
.GLOBAL GND
.end
