magic
tech sky130A
magscale 1 2
timestamp 1725528602
<< pwell >>
rect -1522 -702 1522 702
<< psubdiff >>
rect -1486 632 1486 666
rect -1486 570 -1452 632
rect 1452 570 1486 632
rect -1486 -632 -1452 -570
rect 1452 -632 1486 -570
rect -1486 -666 1486 -632
<< psubdiffcont >>
rect -1486 -570 -1452 570
rect 1452 -570 1486 570
<< xpolycontact >>
rect -1356 104 -1218 536
rect -1356 -536 -1218 -104
rect -1122 104 -984 536
rect -1122 -536 -984 -104
rect -888 104 -750 536
rect -888 -536 -750 -104
rect -654 104 -516 536
rect -654 -536 -516 -104
rect -420 104 -282 536
rect -420 -536 -282 -104
rect -186 104 -48 536
rect -186 -536 -48 -104
rect 48 104 186 536
rect 48 -536 186 -104
rect 282 104 420 536
rect 282 -536 420 -104
rect 516 104 654 536
rect 516 -536 654 -104
rect 750 104 888 536
rect 750 -536 888 -104
rect 984 104 1122 536
rect 984 -536 1122 -104
rect 1218 104 1356 536
rect 1218 -536 1356 -104
<< xpolyres >>
rect -1356 -104 -1218 104
rect -1122 -104 -984 104
rect -888 -104 -750 104
rect -654 -104 -516 104
rect -420 -104 -282 104
rect -186 -104 -48 104
rect 48 -104 186 104
rect 282 -104 420 104
rect 516 -104 654 104
rect 750 -104 888 104
rect 984 -104 1122 104
rect 1218 -104 1356 104
<< locali >>
rect -1486 632 1486 666
rect -1486 570 -1452 632
rect 1452 570 1486 632
rect -1486 -632 -1452 -570
rect 1452 -632 1486 -570
rect -1486 -666 1486 -632
<< viali >>
rect -1340 121 -1234 518
rect -1106 121 -1000 518
rect -872 121 -766 518
rect -638 121 -532 518
rect -404 121 -298 518
rect -170 121 -64 518
rect 64 121 170 518
rect 298 121 404 518
rect 532 121 638 518
rect 766 121 872 518
rect 1000 121 1106 518
rect 1234 121 1340 518
rect -1340 -518 -1234 -121
rect -1106 -518 -1000 -121
rect -872 -518 -766 -121
rect -638 -518 -532 -121
rect -404 -518 -298 -121
rect -170 -518 -64 -121
rect 64 -518 170 -121
rect 298 -518 404 -121
rect 532 -518 638 -121
rect 766 -518 872 -121
rect 1000 -518 1106 -121
rect 1234 -518 1340 -121
<< metal1 >>
rect -1346 518 -1228 530
rect -1346 121 -1340 518
rect -1234 121 -1228 518
rect -1346 109 -1228 121
rect -1112 518 -994 530
rect -1112 121 -1106 518
rect -1000 121 -994 518
rect -1112 109 -994 121
rect -878 518 -760 530
rect -878 121 -872 518
rect -766 121 -760 518
rect -878 109 -760 121
rect -644 518 -526 530
rect -644 121 -638 518
rect -532 121 -526 518
rect -644 109 -526 121
rect -410 518 -292 530
rect -410 121 -404 518
rect -298 121 -292 518
rect -410 109 -292 121
rect -176 518 -58 530
rect -176 121 -170 518
rect -64 121 -58 518
rect -176 109 -58 121
rect 58 518 176 530
rect 58 121 64 518
rect 170 121 176 518
rect 58 109 176 121
rect 292 518 410 530
rect 292 121 298 518
rect 404 121 410 518
rect 292 109 410 121
rect 526 518 644 530
rect 526 121 532 518
rect 638 121 644 518
rect 526 109 644 121
rect 760 518 878 530
rect 760 121 766 518
rect 872 121 878 518
rect 760 109 878 121
rect 994 518 1112 530
rect 994 121 1000 518
rect 1106 121 1112 518
rect 994 109 1112 121
rect 1228 518 1346 530
rect 1228 121 1234 518
rect 1340 121 1346 518
rect 1228 109 1346 121
rect -1346 -121 -1228 -109
rect -1346 -518 -1340 -121
rect -1234 -518 -1228 -121
rect -1346 -530 -1228 -518
rect -1112 -121 -994 -109
rect -1112 -518 -1106 -121
rect -1000 -518 -994 -121
rect -1112 -530 -994 -518
rect -878 -121 -760 -109
rect -878 -518 -872 -121
rect -766 -518 -760 -121
rect -878 -530 -760 -518
rect -644 -121 -526 -109
rect -644 -518 -638 -121
rect -532 -518 -526 -121
rect -644 -530 -526 -518
rect -410 -121 -292 -109
rect -410 -518 -404 -121
rect -298 -518 -292 -121
rect -410 -530 -292 -518
rect -176 -121 -58 -109
rect -176 -518 -170 -121
rect -64 -518 -58 -121
rect -176 -530 -58 -518
rect 58 -121 176 -109
rect 58 -518 64 -121
rect 170 -518 176 -121
rect 58 -530 176 -518
rect 292 -121 410 -109
rect 292 -518 298 -121
rect 404 -518 410 -121
rect 292 -530 410 -518
rect 526 -121 644 -109
rect 526 -518 532 -121
rect 638 -518 644 -121
rect 526 -530 644 -518
rect 760 -121 878 -109
rect 760 -518 766 -121
rect 872 -518 878 -121
rect 760 -530 878 -518
rect 994 -121 1112 -109
rect 994 -518 1000 -121
rect 1106 -518 1112 -121
rect 994 -530 1112 -518
rect 1228 -121 1346 -109
rect 1228 -518 1234 -121
rect 1340 -518 1346 -121
rect 1228 -530 1346 -518
<< properties >>
string FIXED_BBOX -1469 -649 1469 649
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 1.2 m 1 nx 12 wmin 0.690 lmin 0.50 rho 2000 val 4.023k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
