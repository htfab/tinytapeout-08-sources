magic
tech sky130A
magscale 1 2
timestamp 1724945390
<< pwell >>
rect -201 -672 201 672
<< psubdiff >>
rect -165 602 -69 636
rect 69 602 165 636
rect -165 540 -131 602
rect 131 540 165 602
rect -165 -602 -131 -540
rect 131 -602 165 -540
rect -165 -636 -69 -602
rect 69 -636 165 -602
<< psubdiffcont >>
rect -69 602 69 636
rect -165 -540 -131 540
rect 131 -540 165 540
rect -69 -636 69 -602
<< xpolycontact >>
rect -35 74 35 506
rect -35 -506 35 -74
<< xpolyres >>
rect -35 -74 35 74
<< locali >>
rect -165 602 -69 636
rect 69 602 165 636
rect -165 540 -131 602
rect 131 540 165 602
rect -165 -602 -131 -540
rect 131 -602 165 -540
rect -165 -636 -69 -602
rect 69 -636 165 -602
<< viali >>
rect -19 91 19 488
rect -19 -488 19 -91
<< metal1 >>
rect -25 488 25 500
rect -25 91 -19 488
rect 19 91 25 488
rect -25 79 25 91
rect -25 -91 25 -79
rect -25 -488 -19 -91
rect 19 -488 25 -91
rect -25 -500 25 -488
<< properties >>
string FIXED_BBOX -148 -619 148 619
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.9 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 6.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
