magic
tech sky130A
magscale 1 2
timestamp 1725314430
<< pwell >>
rect -2741 -979 2741 979
<< nmoslvt >>
rect -2545 -769 -1745 831
rect -1687 -769 -887 831
rect -829 -769 -29 831
rect 29 -769 829 831
rect 887 -769 1687 831
rect 1745 -769 2545 831
<< ndiff >>
rect -2603 819 -2545 831
rect -2603 -757 -2591 819
rect -2557 -757 -2545 819
rect -2603 -769 -2545 -757
rect -1745 819 -1687 831
rect -1745 -757 -1733 819
rect -1699 -757 -1687 819
rect -1745 -769 -1687 -757
rect -887 819 -829 831
rect -887 -757 -875 819
rect -841 -757 -829 819
rect -887 -769 -829 -757
rect -29 819 29 831
rect -29 -757 -17 819
rect 17 -757 29 819
rect -29 -769 29 -757
rect 829 819 887 831
rect 829 -757 841 819
rect 875 -757 887 819
rect 829 -769 887 -757
rect 1687 819 1745 831
rect 1687 -757 1699 819
rect 1733 -757 1745 819
rect 1687 -769 1745 -757
rect 2545 819 2603 831
rect 2545 -757 2557 819
rect 2591 -757 2603 819
rect 2545 -769 2603 -757
<< ndiffc >>
rect -2591 -757 -2557 819
rect -1733 -757 -1699 819
rect -875 -757 -841 819
rect -17 -757 17 819
rect 841 -757 875 819
rect 1699 -757 1733 819
rect 2557 -757 2591 819
<< psubdiff >>
rect -2705 909 2705 943
rect -2705 847 -2671 909
rect 2671 847 2705 909
rect -2705 -909 -2671 -847
rect 2671 -909 2705 -847
rect -2705 -943 2705 -909
<< psubdiffcont >>
rect -2705 -847 -2671 847
rect 2671 -847 2705 847
<< poly >>
rect -2545 831 -1745 857
rect -1687 831 -887 857
rect -829 831 -29 857
rect 29 831 829 857
rect 887 831 1687 857
rect 1745 831 2545 857
rect -2545 -807 -1745 -769
rect -2545 -841 -2529 -807
rect -1761 -841 -1745 -807
rect -2545 -857 -1745 -841
rect -1687 -807 -887 -769
rect -1687 -841 -1671 -807
rect -903 -841 -887 -807
rect -1687 -857 -887 -841
rect -829 -807 -29 -769
rect -829 -841 -813 -807
rect -45 -841 -29 -807
rect -829 -857 -29 -841
rect 29 -807 829 -769
rect 29 -841 45 -807
rect 813 -841 829 -807
rect 29 -857 829 -841
rect 887 -807 1687 -769
rect 887 -841 903 -807
rect 1671 -841 1687 -807
rect 887 -857 1687 -841
rect 1745 -807 2545 -769
rect 1745 -841 1761 -807
rect 2529 -841 2545 -807
rect 1745 -857 2545 -841
<< polycont >>
rect -2529 -841 -1761 -807
rect -1671 -841 -903 -807
rect -813 -841 -45 -807
rect 45 -841 813 -807
rect 903 -841 1671 -807
rect 1761 -841 2529 -807
<< locali >>
rect -2705 909 2705 943
rect -2705 847 -2671 909
rect 2671 847 2705 909
rect -2591 819 -2557 835
rect -2591 -773 -2557 -757
rect -1733 819 -1699 835
rect -1733 -773 -1699 -757
rect -875 819 -841 835
rect -875 -773 -841 -757
rect -17 819 17 835
rect -17 -773 17 -757
rect 841 819 875 835
rect 841 -773 875 -757
rect 1699 819 1733 835
rect 1699 -773 1733 -757
rect 2557 819 2591 835
rect 2557 -773 2591 -757
rect -2545 -841 -2529 -807
rect -1761 -841 -1745 -807
rect -1687 -841 -1671 -807
rect -903 -841 -887 -807
rect -829 -841 -813 -807
rect -45 -841 -29 -807
rect 29 -841 45 -807
rect 813 -841 829 -807
rect 887 -841 903 -807
rect 1671 -841 1687 -807
rect 1745 -841 1761 -807
rect 2529 -841 2545 -807
rect -2705 -909 -2671 -847
rect 2671 -909 2705 -847
rect -2705 -943 2705 -909
<< viali >>
rect -2591 -740 -2557 -267
rect -1733 329 -1699 802
rect -875 -740 -841 -267
rect -17 329 17 802
rect 841 -740 875 -267
rect 1699 329 1733 802
rect 2557 -740 2591 -267
rect -2529 -841 -1761 -807
rect -1671 -841 -903 -807
rect -813 -841 -45 -807
rect 45 -841 813 -807
rect 903 -841 1671 -807
rect 1761 -841 2529 -807
<< metal1 >>
rect -1739 802 -1693 814
rect -1739 329 -1733 802
rect -1699 329 -1693 802
rect -1739 317 -1693 329
rect -23 802 23 814
rect -23 329 -17 802
rect 17 329 23 802
rect -23 317 23 329
rect 1693 802 1739 814
rect 1693 329 1699 802
rect 1733 329 1739 802
rect 1693 317 1739 329
rect -2597 -267 -2551 -255
rect -2597 -740 -2591 -267
rect -2557 -740 -2551 -267
rect -2597 -752 -2551 -740
rect -881 -267 -835 -255
rect -881 -740 -875 -267
rect -841 -740 -835 -267
rect -881 -752 -835 -740
rect 835 -267 881 -255
rect 835 -740 841 -267
rect 875 -740 881 -267
rect 835 -752 881 -740
rect 2551 -267 2597 -255
rect 2551 -740 2557 -267
rect 2591 -740 2597 -267
rect 2551 -752 2597 -740
rect -2541 -807 -1749 -801
rect -2541 -841 -2529 -807
rect -1761 -841 -1749 -807
rect -2541 -847 -1749 -841
rect -1683 -807 -891 -801
rect -1683 -841 -1671 -807
rect -903 -841 -891 -807
rect -1683 -847 -891 -841
rect -825 -807 -33 -801
rect -825 -841 -813 -807
rect -45 -841 -33 -807
rect -825 -847 -33 -841
rect 33 -807 825 -801
rect 33 -841 45 -807
rect 813 -841 825 -807
rect 33 -847 825 -841
rect 891 -807 1683 -801
rect 891 -841 903 -807
rect 1671 -841 1683 -807
rect 891 -847 1683 -841
rect 1749 -807 2541 -801
rect 1749 -841 1761 -807
rect 2529 -841 2541 -807
rect 1749 -847 2541 -841
<< properties >>
string FIXED_BBOX -2688 -926 2688 926
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8 l 4 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -30 viadrn +30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
