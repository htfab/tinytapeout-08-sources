magic
tech sky130A
magscale 1 2
timestamp 1725467640
<< nwell >>
rect -2804 -199 -1202 -195
rect -2908 -1599 -1202 -199
rect -2804 -1602 -1202 -1599
<< psubdiff >>
rect 6539 -580 6738 -463
rect 6539 -1212 6603 -580
rect 6675 -1212 6738 -580
rect 6539 -1393 6738 -1212
<< nsubdiff >>
rect -2783 -433 -2621 -393
rect -2783 -1338 -2746 -433
rect -2661 -1338 -2621 -433
rect -2783 -1397 -2621 -1338
rect -1401 -429 -1239 -397
rect -1401 -1334 -1356 -429
rect -1271 -1334 -1239 -429
rect -1401 -1401 -1239 -1334
<< psubdiffcont >>
rect 6603 -1212 6675 -580
<< nsubdiffcont >>
rect -2746 -1338 -2661 -433
rect -1356 -1334 -1271 -429
<< locali >>
rect -2760 -433 -2647 -411
rect -2760 -1338 -2746 -433
rect -2661 -537 -2647 -433
rect -2651 -789 -2647 -537
rect -2661 -1338 -2647 -789
rect -2760 -1388 -2647 -1338
rect -1378 -429 -1265 -411
rect -1378 -546 -1356 -429
rect -1271 -546 -1265 -429
rect -1378 -798 -1365 -546
rect -1270 -798 -1265 -546
rect -1378 -1334 -1356 -798
rect -1271 -1334 -1265 -798
rect 6576 -580 6711 -526
rect 6576 -722 6603 -580
rect 6675 -722 6711 -580
rect 6576 -865 6584 -722
rect 6576 -1212 6603 -865
rect 6675 -1212 6711 -865
rect 6576 -1312 6711 -1212
rect -1378 -1388 -1265 -1334
<< viali >>
rect -2746 -789 -2661 -537
rect -2661 -789 -2651 -537
rect -1365 -798 -1356 -546
rect -1356 -798 -1271 -546
rect -1271 -798 -1270 -546
rect 6584 -865 6603 -722
rect 6603 -865 6675 -722
rect 6675 -865 6727 -722
<< metal1 >>
rect -2509 -405 -1529 -395
rect -2759 -804 -2749 -428
rect -2643 -546 -2633 -428
rect -2509 -507 -2322 -405
rect -2239 -507 -1529 -405
rect -2509 -517 -1529 -507
rect -1381 -546 -1371 -423
rect -2643 -799 -1371 -546
rect -1265 -799 -1255 -423
rect 6193 -506 6541 -503
rect -2643 -802 -1264 -799
rect -2643 -804 -2633 -802
rect -1371 -810 -1264 -802
rect -621 -830 6541 -506
rect -621 -831 6321 -830
rect 6420 -965 6541 -830
rect 6572 -722 7170 -716
rect 6572 -865 6584 -722
rect 6727 -865 7170 -722
rect 6572 -871 7170 -865
rect 5380 -1039 5386 -1034
rect 245 -1043 2006 -1039
rect 3694 -1043 5386 -1039
rect -2328 -1055 -2228 -1048
rect -2332 -1319 -2322 -1055
rect -2239 -1319 -2228 -1055
rect -2328 -1666 -2228 -1319
rect -1813 -1467 -1713 -1048
rect 234 -1143 240 -1043
rect 340 -1052 2006 -1043
rect 340 -1143 1947 -1052
rect 245 -1152 1947 -1143
rect 2047 -1152 2053 -1052
rect 3656 -1143 3662 -1043
rect 3762 -1134 5386 -1043
rect 5486 -1134 5492 -1034
rect 6420 -1086 7005 -965
rect 3762 -1143 5455 -1134
rect 7276 -1140 7332 -959
rect 245 -1301 2006 -1152
rect 3694 -1301 5455 -1143
rect 6858 -1199 7332 -1140
rect -558 -1539 2818 -1332
rect 2890 -1541 6266 -1334
rect -1813 -1573 -1713 -1567
rect 240 -1666 340 -1660
rect -2328 -1766 240 -1666
rect 340 -1766 1947 -1666
rect 2047 -1766 2053 -1666
rect 240 -1772 340 -1766
<< via1 >>
rect -2749 -537 -2643 -428
rect -2749 -789 -2746 -537
rect -2746 -789 -2651 -537
rect -2651 -789 -2643 -537
rect -2322 -507 -2239 -405
rect -1371 -546 -1265 -423
rect -2749 -804 -2643 -789
rect -1371 -798 -1365 -546
rect -1365 -798 -1270 -546
rect -1270 -798 -1265 -546
rect -1371 -799 -1265 -798
rect -2322 -1319 -2239 -1055
rect 240 -1143 340 -1043
rect 1947 -1152 2047 -1052
rect 3662 -1143 3762 -1043
rect 5386 -1134 5486 -1034
rect -1813 -1567 -1713 -1467
rect 240 -1766 340 -1666
rect 1947 -1766 2047 -1666
<< metal2 >>
rect -2322 -398 -2239 -395
rect -2332 -405 -2225 -398
rect -2749 -428 -2643 -418
rect -2749 -814 -2643 -804
rect -2332 -507 -2322 -405
rect -2239 -507 -2225 -405
rect -2332 -1055 -2225 -507
rect -1371 -423 -1265 -413
rect -1371 -809 -1265 -799
rect 5386 -1034 5486 -1028
rect -2332 -1319 -2322 -1055
rect -2239 -1319 -2225 -1055
rect -2332 -1333 -2225 -1319
rect 240 -1043 340 -1037
rect 3662 -1043 3762 -1037
rect -1819 -1567 -1813 -1467
rect -1713 -1567 -1707 -1467
rect -1813 -1828 -1713 -1567
rect 240 -1666 340 -1143
rect 1947 -1052 2047 -1046
rect 1947 -1666 2047 -1152
rect 234 -1766 240 -1666
rect 340 -1766 346 -1666
rect 1947 -1772 2047 -1766
rect 3662 -1828 3762 -1143
rect 5386 -1828 5486 -1134
rect -1813 -1928 5486 -1828
<< via2 >>
rect -2749 -804 -2643 -428
rect -1371 -799 -1265 -423
<< metal3 >>
rect -2759 73 -1253 203
rect -2759 -428 -2629 73
rect -2759 -804 -2749 -428
rect -2643 -794 -2629 -428
rect -1383 -423 -1253 73
rect -2643 -804 -2633 -794
rect -1383 -799 -1371 -423
rect -1265 -799 -1253 -423
rect -1383 -801 -1253 -799
rect -1381 -804 -1255 -801
rect -2759 -809 -2633 -804
use sky130_fd_pr__nfet_01v8_lvt_DG3K4W  sky130_fd_pr__nfet_01v8_lvt_DG3K4W_0
timestamp 1725467580
transform 1 0 7066 0 1 -943
box -266 -257 266 257
use sky130_fd_pr__nfet_01v8_lvt_LJJETC  sky130_fd_pr__nfet_01v8_lvt_LJJETC_0
timestamp 1725467580
transform 1 0 2858 0 1 -945
box -3461 -457 3461 457
use sky130_fd_pr__pfet_01v8_lvt_EBPRJ2  sky130_fd_pr__pfet_01v8_lvt_EBPRJ2_0
timestamp 1725467580
transform 1 0 -2019 0 1 -904
box -581 -498 581 464
<< labels >>
flabel metal3 -2219 97 -2036 184 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 -451 -1531 -253 -1425 0 FreeSans 160 0 0 0 PLUS
port 5 nsew
flabel metal1 3052 -1522 3293 -1420 0 FreeSans 160 0 0 0 MINUS
port 4 nsew
flabel metal1 6743 -859 6798 -723 0 FreeSans 160 90 0 0 VSS
port 2 nsew
flabel metal1 7279 -1192 7320 -1135 0 FreeSans 80 90 0 0 in
port 3 nsew
flabel metal2 4469 -1909 4604 -1836 0 FreeSans 160 0 0 0 opout
port 6 nsew
<< end >>
