magic
tech sky130A
magscale 1 2
timestamp 1725569918
<< pwell >>
rect -625 -410 625 410
<< nmos >>
rect -429 -200 -29 200
rect 29 -200 429 200
<< ndiff >>
rect -487 188 -429 200
rect -487 -188 -475 188
rect -441 -188 -429 188
rect -487 -200 -429 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 429 188 487 200
rect 429 -188 441 188
rect 475 -188 487 188
rect 429 -200 487 -188
<< ndiffc >>
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
<< psubdiff >>
rect -589 340 -493 374
rect 493 340 589 374
rect -589 278 -555 340
rect 555 278 589 340
rect -589 -340 -555 -278
rect 555 -340 589 -278
rect -589 -374 -493 -340
rect 493 -374 589 -340
<< psubdiffcont >>
rect -493 340 493 374
rect -589 -278 -555 278
rect 555 -278 589 278
rect -493 -374 493 -340
<< poly >>
rect -429 272 -29 288
rect -429 238 -413 272
rect -45 238 -29 272
rect -429 200 -29 238
rect 29 272 429 288
rect 29 238 45 272
rect 413 238 429 272
rect 29 200 429 238
rect -429 -238 -29 -200
rect -429 -272 -413 -238
rect -45 -272 -29 -238
rect -429 -288 -29 -272
rect 29 -238 429 -200
rect 29 -272 45 -238
rect 413 -272 429 -238
rect 29 -288 429 -272
<< polycont >>
rect -413 238 -45 272
rect 45 238 413 272
rect -413 -272 -45 -238
rect 45 -272 413 -238
<< locali >>
rect -589 340 -493 374
rect 493 340 589 374
rect -589 278 -555 340
rect 555 278 589 340
rect -429 238 -413 272
rect -45 238 -29 272
rect 29 238 45 272
rect 413 238 429 272
rect -475 188 -441 204
rect -475 -204 -441 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 441 188 475 204
rect 441 -204 475 -188
rect -429 -272 -413 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 413 -272 429 -238
rect -589 -340 -555 -278
rect 555 -340 589 -278
rect -589 -374 -493 -340
rect 493 -374 589 -340
<< viali >>
rect -413 238 -45 272
rect 45 238 413 272
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect -413 -272 -45 -238
rect 45 -272 413 -238
<< metal1 >>
rect -425 272 -33 278
rect -425 238 -413 272
rect -45 238 -33 272
rect -425 232 -33 238
rect 33 272 425 278
rect 33 238 45 272
rect 413 238 425 272
rect 33 232 425 238
rect -481 188 -435 200
rect -481 -188 -475 188
rect -441 -188 -435 188
rect -481 -200 -435 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 435 188 481 200
rect 435 -188 441 188
rect 475 -188 481 188
rect 435 -200 481 -188
rect -425 -238 -33 -232
rect -425 -272 -413 -238
rect -45 -272 -33 -238
rect -425 -278 -33 -272
rect 33 -238 425 -232
rect 33 -272 45 -238
rect 413 -272 425 -238
rect 33 -278 425 -272
<< properties >>
string FIXED_BBOX -572 -357 572 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 2.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
