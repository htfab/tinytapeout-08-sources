** sch_path: /home/ttuser/test0/tt08-bgr/xschem/core_prel.sch
.subckt core_prel VDD Vbgr VSS
*.PININFO VDD:I VSS:I Vbgr:O
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40  m=1
XQ2 VSS VSS net1 sky130_fd_pr__pnp_05v5_W3p40L3p40   m=29
XM1 MINUS opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM2 PLUS opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM3 Vbgr opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XM4 opout MINUS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 m=1
XM5 Gcm1 PLUS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 m=1
XM6 opout Gcm1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
XM10 Sop Gcm2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 m=1
XM9 Gcm2 Gcm2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 m=1
XM7 Gcm1 Gcm1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
XM8 Gcm2 opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 m=1
XR19 net1 PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.05 mult=1 m=1
XR3 VSS MINUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6 mult=1 m=1
XR4 VSS Vbgr VSS sky130_fd_pr__res_xhigh_po_0p69 L=12.6 mult=1 m=1
XM12 VSS Vbgr opout opout sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=4
XR2 VSS PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6 mult=1 m=1
XR1 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XR5 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
XR6 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p69 L=1.26 mult=1 m=1
XM17 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=5 nf=1 m=1
XM18 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 m=1
XM19 Gcm2 VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 m=1
XR7 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p69 L=1.26 mult=1 m=1
XM20 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=1
XR8 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.05 mult=1 m=1
XR9 VSS VSS VSS sky130_fd_pr__res_xhigh_po_0p35 L=1.05 mult=1 m=1
XM21 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=1
XM11 VSS VSS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=8 nf=1 m=1
XM13 VSS VSS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=8 nf=1 m=1
XM14 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=5 nf=1 m=1
XM15 opout VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XM16 opout VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
.ends
.end
