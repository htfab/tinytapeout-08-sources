magic
tech sky130A
magscale 1 2
timestamp 1725572295
<< locali >>
rect 520 -80 3230 200
rect 520 -810 730 -80
rect 1900 -810 1970 -80
rect 3140 -810 3230 -80
rect 520 -910 3230 -810
rect 520 -1000 900 -910
rect 3160 -1000 3230 -910
rect 520 -1060 3230 -1000
rect 3300 150 4290 200
rect 3300 -1010 3650 150
rect 4010 -830 4150 150
rect 4240 -830 4290 150
rect 4010 -1010 4290 -830
rect 3300 -1060 4290 -1010
<< viali >>
rect 900 -1000 3160 -910
rect 4150 -830 4240 150
<< metal1 >>
rect 520 180 3230 200
rect 520 10 1280 180
rect 1350 10 3230 180
rect 520 0 3230 10
rect 3300 70 3500 200
rect 4090 150 4290 200
rect 3300 0 3870 70
rect 790 -860 840 -240
rect 1020 -720 1150 0
rect 1270 -250 1360 -240
rect 1270 -630 1280 -250
rect 1350 -630 1360 -250
rect 1270 -640 1360 -630
rect 1480 -710 1610 0
rect 1790 -860 1840 -240
rect 2030 -860 2080 -240
rect 2280 -720 2410 0
rect 2510 -260 2600 -250
rect 2510 -640 2520 -260
rect 2590 -640 2600 -260
rect 2510 -650 2600 -640
rect 2730 -710 2860 0
rect 3030 -860 3080 -240
rect 3300 -260 3500 0
rect 3300 -640 3360 -260
rect 3430 -410 3500 -260
rect 4090 -410 4150 150
rect 3430 -480 3800 -410
rect 3860 -480 4150 -410
rect 3430 -640 3500 -480
rect 3300 -860 3500 -640
rect 4090 -830 4150 -480
rect 4240 -830 4290 150
rect 520 -910 3230 -860
rect 520 -1000 900 -910
rect 3160 -1000 3230 -910
rect 520 -1060 3230 -1000
rect 3300 -930 3870 -860
rect 3300 -1060 3500 -930
rect 4090 -1060 4290 -830
<< via1 >>
rect 1280 10 1350 180
rect 1280 -630 1350 -250
rect 2520 -640 2590 -260
rect 3360 -640 3430 -260
<< metal2 >>
rect 1270 180 1360 190
rect 1270 10 1280 180
rect 1350 10 1360 180
rect 1270 -250 1360 10
rect 1270 -630 1280 -250
rect 1350 -630 1360 -250
rect 1270 -640 1360 -630
rect 2510 -260 2600 -250
rect 2510 -640 2520 -260
rect 2590 -410 2600 -260
rect 3350 -260 3440 -250
rect 3350 -410 3360 -260
rect 2590 -480 3360 -410
rect 2590 -640 2600 -480
rect 2510 -650 2600 -640
rect 3350 -640 3360 -480
rect 3430 -640 3440 -260
rect 3350 -650 3440 -640
use sky130_fd_pr__nfet_01v8_XVWV9B  XM1
timestamp 1725569918
transform 1 0 1315 0 1 -440
box -625 -410 625 410
use sky130_fd_pr__nfet_01v8_XVWV9B  XM2
timestamp 1725569918
transform 1 0 2555 0 1 -450
box -625 -410 625 410
use sky130_fd_pr__pfet_01v8_NDBSV3  XM3
timestamp 1725569918
transform 1 0 3831 0 1 -431
box -221 -619 221 619
<< labels >>
flabel metal1 520 -1060 720 -860 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 520 0 720 200 0 FreeSans 256 0 0 0 Icont
port 2 nsew
flabel metal1 3300 -1060 3500 -860 0 FreeSans 256 0 0 0 Vb
port 3 nsew
flabel metal1 4090 -1060 4290 -860 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
