magic
tech sky130A
magscale 1 2
timestamp 1723635744
<< metal3 >>
rect -436 40852 436 40880
rect -436 40328 352 40852
rect 416 40328 436 40852
rect -436 40300 436 40328
rect -436 40032 436 40060
rect -436 39508 352 40032
rect 416 39508 436 40032
rect -436 39480 436 39508
rect -436 39212 436 39240
rect -436 38688 352 39212
rect 416 38688 436 39212
rect -436 38660 436 38688
rect -436 38392 436 38420
rect -436 37868 352 38392
rect 416 37868 436 38392
rect -436 37840 436 37868
rect -436 37572 436 37600
rect -436 37048 352 37572
rect 416 37048 436 37572
rect -436 37020 436 37048
rect -436 36752 436 36780
rect -436 36228 352 36752
rect 416 36228 436 36752
rect -436 36200 436 36228
rect -436 35932 436 35960
rect -436 35408 352 35932
rect 416 35408 436 35932
rect -436 35380 436 35408
rect -436 35112 436 35140
rect -436 34588 352 35112
rect 416 34588 436 35112
rect -436 34560 436 34588
rect -436 34292 436 34320
rect -436 33768 352 34292
rect 416 33768 436 34292
rect -436 33740 436 33768
rect -436 33472 436 33500
rect -436 32948 352 33472
rect 416 32948 436 33472
rect -436 32920 436 32948
rect -436 32652 436 32680
rect -436 32128 352 32652
rect 416 32128 436 32652
rect -436 32100 436 32128
rect -436 31832 436 31860
rect -436 31308 352 31832
rect 416 31308 436 31832
rect -436 31280 436 31308
rect -436 31012 436 31040
rect -436 30488 352 31012
rect 416 30488 436 31012
rect -436 30460 436 30488
rect -436 30192 436 30220
rect -436 29668 352 30192
rect 416 29668 436 30192
rect -436 29640 436 29668
rect -436 29372 436 29400
rect -436 28848 352 29372
rect 416 28848 436 29372
rect -436 28820 436 28848
rect -436 28552 436 28580
rect -436 28028 352 28552
rect 416 28028 436 28552
rect -436 28000 436 28028
rect -436 27732 436 27760
rect -436 27208 352 27732
rect 416 27208 436 27732
rect -436 27180 436 27208
rect -436 26912 436 26940
rect -436 26388 352 26912
rect 416 26388 436 26912
rect -436 26360 436 26388
rect -436 26092 436 26120
rect -436 25568 352 26092
rect 416 25568 436 26092
rect -436 25540 436 25568
rect -436 25272 436 25300
rect -436 24748 352 25272
rect 416 24748 436 25272
rect -436 24720 436 24748
rect -436 24452 436 24480
rect -436 23928 352 24452
rect 416 23928 436 24452
rect -436 23900 436 23928
rect -436 23632 436 23660
rect -436 23108 352 23632
rect 416 23108 436 23632
rect -436 23080 436 23108
rect -436 22812 436 22840
rect -436 22288 352 22812
rect 416 22288 436 22812
rect -436 22260 436 22288
rect -436 21992 436 22020
rect -436 21468 352 21992
rect 416 21468 436 21992
rect -436 21440 436 21468
rect -436 21172 436 21200
rect -436 20648 352 21172
rect 416 20648 436 21172
rect -436 20620 436 20648
rect -436 20352 436 20380
rect -436 19828 352 20352
rect 416 19828 436 20352
rect -436 19800 436 19828
rect -436 19532 436 19560
rect -436 19008 352 19532
rect 416 19008 436 19532
rect -436 18980 436 19008
rect -436 18712 436 18740
rect -436 18188 352 18712
rect 416 18188 436 18712
rect -436 18160 436 18188
rect -436 17892 436 17920
rect -436 17368 352 17892
rect 416 17368 436 17892
rect -436 17340 436 17368
rect -436 17072 436 17100
rect -436 16548 352 17072
rect 416 16548 436 17072
rect -436 16520 436 16548
rect -436 16252 436 16280
rect -436 15728 352 16252
rect 416 15728 436 16252
rect -436 15700 436 15728
rect -436 15432 436 15460
rect -436 14908 352 15432
rect 416 14908 436 15432
rect -436 14880 436 14908
rect -436 14612 436 14640
rect -436 14088 352 14612
rect 416 14088 436 14612
rect -436 14060 436 14088
rect -436 13792 436 13820
rect -436 13268 352 13792
rect 416 13268 436 13792
rect -436 13240 436 13268
rect -436 12972 436 13000
rect -436 12448 352 12972
rect 416 12448 436 12972
rect -436 12420 436 12448
rect -436 12152 436 12180
rect -436 11628 352 12152
rect 416 11628 436 12152
rect -436 11600 436 11628
rect -436 11332 436 11360
rect -436 10808 352 11332
rect 416 10808 436 11332
rect -436 10780 436 10808
rect -436 10512 436 10540
rect -436 9988 352 10512
rect 416 9988 436 10512
rect -436 9960 436 9988
rect -436 9692 436 9720
rect -436 9168 352 9692
rect 416 9168 436 9692
rect -436 9140 436 9168
rect -436 8872 436 8900
rect -436 8348 352 8872
rect 416 8348 436 8872
rect -436 8320 436 8348
rect -436 8052 436 8080
rect -436 7528 352 8052
rect 416 7528 436 8052
rect -436 7500 436 7528
rect -436 7232 436 7260
rect -436 6708 352 7232
rect 416 6708 436 7232
rect -436 6680 436 6708
rect -436 6412 436 6440
rect -436 5888 352 6412
rect 416 5888 436 6412
rect -436 5860 436 5888
rect -436 5592 436 5620
rect -436 5068 352 5592
rect 416 5068 436 5592
rect -436 5040 436 5068
rect -436 4772 436 4800
rect -436 4248 352 4772
rect 416 4248 436 4772
rect -436 4220 436 4248
rect -436 3952 436 3980
rect -436 3428 352 3952
rect 416 3428 436 3952
rect -436 3400 436 3428
rect -436 3132 436 3160
rect -436 2608 352 3132
rect 416 2608 436 3132
rect -436 2580 436 2608
rect -436 2312 436 2340
rect -436 1788 352 2312
rect 416 1788 436 2312
rect -436 1760 436 1788
rect -436 1492 436 1520
rect -436 968 352 1492
rect 416 968 436 1492
rect -436 940 436 968
rect -436 672 436 700
rect -436 148 352 672
rect 416 148 436 672
rect -436 120 436 148
rect -436 -148 436 -120
rect -436 -672 352 -148
rect 416 -672 436 -148
rect -436 -700 436 -672
rect -436 -968 436 -940
rect -436 -1492 352 -968
rect 416 -1492 436 -968
rect -436 -1520 436 -1492
rect -436 -1788 436 -1760
rect -436 -2312 352 -1788
rect 416 -2312 436 -1788
rect -436 -2340 436 -2312
rect -436 -2608 436 -2580
rect -436 -3132 352 -2608
rect 416 -3132 436 -2608
rect -436 -3160 436 -3132
rect -436 -3428 436 -3400
rect -436 -3952 352 -3428
rect 416 -3952 436 -3428
rect -436 -3980 436 -3952
rect -436 -4248 436 -4220
rect -436 -4772 352 -4248
rect 416 -4772 436 -4248
rect -436 -4800 436 -4772
rect -436 -5068 436 -5040
rect -436 -5592 352 -5068
rect 416 -5592 436 -5068
rect -436 -5620 436 -5592
rect -436 -5888 436 -5860
rect -436 -6412 352 -5888
rect 416 -6412 436 -5888
rect -436 -6440 436 -6412
rect -436 -6708 436 -6680
rect -436 -7232 352 -6708
rect 416 -7232 436 -6708
rect -436 -7260 436 -7232
rect -436 -7528 436 -7500
rect -436 -8052 352 -7528
rect 416 -8052 436 -7528
rect -436 -8080 436 -8052
rect -436 -8348 436 -8320
rect -436 -8872 352 -8348
rect 416 -8872 436 -8348
rect -436 -8900 436 -8872
rect -436 -9168 436 -9140
rect -436 -9692 352 -9168
rect 416 -9692 436 -9168
rect -436 -9720 436 -9692
rect -436 -9988 436 -9960
rect -436 -10512 352 -9988
rect 416 -10512 436 -9988
rect -436 -10540 436 -10512
rect -436 -10808 436 -10780
rect -436 -11332 352 -10808
rect 416 -11332 436 -10808
rect -436 -11360 436 -11332
rect -436 -11628 436 -11600
rect -436 -12152 352 -11628
rect 416 -12152 436 -11628
rect -436 -12180 436 -12152
rect -436 -12448 436 -12420
rect -436 -12972 352 -12448
rect 416 -12972 436 -12448
rect -436 -13000 436 -12972
rect -436 -13268 436 -13240
rect -436 -13792 352 -13268
rect 416 -13792 436 -13268
rect -436 -13820 436 -13792
rect -436 -14088 436 -14060
rect -436 -14612 352 -14088
rect 416 -14612 436 -14088
rect -436 -14640 436 -14612
rect -436 -14908 436 -14880
rect -436 -15432 352 -14908
rect 416 -15432 436 -14908
rect -436 -15460 436 -15432
rect -436 -15728 436 -15700
rect -436 -16252 352 -15728
rect 416 -16252 436 -15728
rect -436 -16280 436 -16252
rect -436 -16548 436 -16520
rect -436 -17072 352 -16548
rect 416 -17072 436 -16548
rect -436 -17100 436 -17072
rect -436 -17368 436 -17340
rect -436 -17892 352 -17368
rect 416 -17892 436 -17368
rect -436 -17920 436 -17892
rect -436 -18188 436 -18160
rect -436 -18712 352 -18188
rect 416 -18712 436 -18188
rect -436 -18740 436 -18712
rect -436 -19008 436 -18980
rect -436 -19532 352 -19008
rect 416 -19532 436 -19008
rect -436 -19560 436 -19532
rect -436 -19828 436 -19800
rect -436 -20352 352 -19828
rect 416 -20352 436 -19828
rect -436 -20380 436 -20352
rect -436 -20648 436 -20620
rect -436 -21172 352 -20648
rect 416 -21172 436 -20648
rect -436 -21200 436 -21172
rect -436 -21468 436 -21440
rect -436 -21992 352 -21468
rect 416 -21992 436 -21468
rect -436 -22020 436 -21992
rect -436 -22288 436 -22260
rect -436 -22812 352 -22288
rect 416 -22812 436 -22288
rect -436 -22840 436 -22812
rect -436 -23108 436 -23080
rect -436 -23632 352 -23108
rect 416 -23632 436 -23108
rect -436 -23660 436 -23632
rect -436 -23928 436 -23900
rect -436 -24452 352 -23928
rect 416 -24452 436 -23928
rect -436 -24480 436 -24452
rect -436 -24748 436 -24720
rect -436 -25272 352 -24748
rect 416 -25272 436 -24748
rect -436 -25300 436 -25272
rect -436 -25568 436 -25540
rect -436 -26092 352 -25568
rect 416 -26092 436 -25568
rect -436 -26120 436 -26092
rect -436 -26388 436 -26360
rect -436 -26912 352 -26388
rect 416 -26912 436 -26388
rect -436 -26940 436 -26912
rect -436 -27208 436 -27180
rect -436 -27732 352 -27208
rect 416 -27732 436 -27208
rect -436 -27760 436 -27732
rect -436 -28028 436 -28000
rect -436 -28552 352 -28028
rect 416 -28552 436 -28028
rect -436 -28580 436 -28552
rect -436 -28848 436 -28820
rect -436 -29372 352 -28848
rect 416 -29372 436 -28848
rect -436 -29400 436 -29372
rect -436 -29668 436 -29640
rect -436 -30192 352 -29668
rect 416 -30192 436 -29668
rect -436 -30220 436 -30192
rect -436 -30488 436 -30460
rect -436 -31012 352 -30488
rect 416 -31012 436 -30488
rect -436 -31040 436 -31012
rect -436 -31308 436 -31280
rect -436 -31832 352 -31308
rect 416 -31832 436 -31308
rect -436 -31860 436 -31832
rect -436 -32128 436 -32100
rect -436 -32652 352 -32128
rect 416 -32652 436 -32128
rect -436 -32680 436 -32652
rect -436 -32948 436 -32920
rect -436 -33472 352 -32948
rect 416 -33472 436 -32948
rect -436 -33500 436 -33472
rect -436 -33768 436 -33740
rect -436 -34292 352 -33768
rect 416 -34292 436 -33768
rect -436 -34320 436 -34292
rect -436 -34588 436 -34560
rect -436 -35112 352 -34588
rect 416 -35112 436 -34588
rect -436 -35140 436 -35112
rect -436 -35408 436 -35380
rect -436 -35932 352 -35408
rect 416 -35932 436 -35408
rect -436 -35960 436 -35932
rect -436 -36228 436 -36200
rect -436 -36752 352 -36228
rect 416 -36752 436 -36228
rect -436 -36780 436 -36752
rect -436 -37048 436 -37020
rect -436 -37572 352 -37048
rect 416 -37572 436 -37048
rect -436 -37600 436 -37572
rect -436 -37868 436 -37840
rect -436 -38392 352 -37868
rect 416 -38392 436 -37868
rect -436 -38420 436 -38392
rect -436 -38688 436 -38660
rect -436 -39212 352 -38688
rect 416 -39212 436 -38688
rect -436 -39240 436 -39212
rect -436 -39508 436 -39480
rect -436 -40032 352 -39508
rect 416 -40032 436 -39508
rect -436 -40060 436 -40032
rect -436 -40328 436 -40300
rect -436 -40852 352 -40328
rect 416 -40852 436 -40328
rect -436 -40880 436 -40852
<< via3 >>
rect 352 40328 416 40852
rect 352 39508 416 40032
rect 352 38688 416 39212
rect 352 37868 416 38392
rect 352 37048 416 37572
rect 352 36228 416 36752
rect 352 35408 416 35932
rect 352 34588 416 35112
rect 352 33768 416 34292
rect 352 32948 416 33472
rect 352 32128 416 32652
rect 352 31308 416 31832
rect 352 30488 416 31012
rect 352 29668 416 30192
rect 352 28848 416 29372
rect 352 28028 416 28552
rect 352 27208 416 27732
rect 352 26388 416 26912
rect 352 25568 416 26092
rect 352 24748 416 25272
rect 352 23928 416 24452
rect 352 23108 416 23632
rect 352 22288 416 22812
rect 352 21468 416 21992
rect 352 20648 416 21172
rect 352 19828 416 20352
rect 352 19008 416 19532
rect 352 18188 416 18712
rect 352 17368 416 17892
rect 352 16548 416 17072
rect 352 15728 416 16252
rect 352 14908 416 15432
rect 352 14088 416 14612
rect 352 13268 416 13792
rect 352 12448 416 12972
rect 352 11628 416 12152
rect 352 10808 416 11332
rect 352 9988 416 10512
rect 352 9168 416 9692
rect 352 8348 416 8872
rect 352 7528 416 8052
rect 352 6708 416 7232
rect 352 5888 416 6412
rect 352 5068 416 5592
rect 352 4248 416 4772
rect 352 3428 416 3952
rect 352 2608 416 3132
rect 352 1788 416 2312
rect 352 968 416 1492
rect 352 148 416 672
rect 352 -672 416 -148
rect 352 -1492 416 -968
rect 352 -2312 416 -1788
rect 352 -3132 416 -2608
rect 352 -3952 416 -3428
rect 352 -4772 416 -4248
rect 352 -5592 416 -5068
rect 352 -6412 416 -5888
rect 352 -7232 416 -6708
rect 352 -8052 416 -7528
rect 352 -8872 416 -8348
rect 352 -9692 416 -9168
rect 352 -10512 416 -9988
rect 352 -11332 416 -10808
rect 352 -12152 416 -11628
rect 352 -12972 416 -12448
rect 352 -13792 416 -13268
rect 352 -14612 416 -14088
rect 352 -15432 416 -14908
rect 352 -16252 416 -15728
rect 352 -17072 416 -16548
rect 352 -17892 416 -17368
rect 352 -18712 416 -18188
rect 352 -19532 416 -19008
rect 352 -20352 416 -19828
rect 352 -21172 416 -20648
rect 352 -21992 416 -21468
rect 352 -22812 416 -22288
rect 352 -23632 416 -23108
rect 352 -24452 416 -23928
rect 352 -25272 416 -24748
rect 352 -26092 416 -25568
rect 352 -26912 416 -26388
rect 352 -27732 416 -27208
rect 352 -28552 416 -28028
rect 352 -29372 416 -28848
rect 352 -30192 416 -29668
rect 352 -31012 416 -30488
rect 352 -31832 416 -31308
rect 352 -32652 416 -32128
rect 352 -33472 416 -32948
rect 352 -34292 416 -33768
rect 352 -35112 416 -34588
rect 352 -35932 416 -35408
rect 352 -36752 416 -36228
rect 352 -37572 416 -37048
rect 352 -38392 416 -37868
rect 352 -39212 416 -38688
rect 352 -40032 416 -39508
rect 352 -40852 416 -40328
<< mimcap >>
rect -396 40800 104 40840
rect -396 40380 -356 40800
rect 64 40380 104 40800
rect -396 40340 104 40380
rect -396 39980 104 40020
rect -396 39560 -356 39980
rect 64 39560 104 39980
rect -396 39520 104 39560
rect -396 39160 104 39200
rect -396 38740 -356 39160
rect 64 38740 104 39160
rect -396 38700 104 38740
rect -396 38340 104 38380
rect -396 37920 -356 38340
rect 64 37920 104 38340
rect -396 37880 104 37920
rect -396 37520 104 37560
rect -396 37100 -356 37520
rect 64 37100 104 37520
rect -396 37060 104 37100
rect -396 36700 104 36740
rect -396 36280 -356 36700
rect 64 36280 104 36700
rect -396 36240 104 36280
rect -396 35880 104 35920
rect -396 35460 -356 35880
rect 64 35460 104 35880
rect -396 35420 104 35460
rect -396 35060 104 35100
rect -396 34640 -356 35060
rect 64 34640 104 35060
rect -396 34600 104 34640
rect -396 34240 104 34280
rect -396 33820 -356 34240
rect 64 33820 104 34240
rect -396 33780 104 33820
rect -396 33420 104 33460
rect -396 33000 -356 33420
rect 64 33000 104 33420
rect -396 32960 104 33000
rect -396 32600 104 32640
rect -396 32180 -356 32600
rect 64 32180 104 32600
rect -396 32140 104 32180
rect -396 31780 104 31820
rect -396 31360 -356 31780
rect 64 31360 104 31780
rect -396 31320 104 31360
rect -396 30960 104 31000
rect -396 30540 -356 30960
rect 64 30540 104 30960
rect -396 30500 104 30540
rect -396 30140 104 30180
rect -396 29720 -356 30140
rect 64 29720 104 30140
rect -396 29680 104 29720
rect -396 29320 104 29360
rect -396 28900 -356 29320
rect 64 28900 104 29320
rect -396 28860 104 28900
rect -396 28500 104 28540
rect -396 28080 -356 28500
rect 64 28080 104 28500
rect -396 28040 104 28080
rect -396 27680 104 27720
rect -396 27260 -356 27680
rect 64 27260 104 27680
rect -396 27220 104 27260
rect -396 26860 104 26900
rect -396 26440 -356 26860
rect 64 26440 104 26860
rect -396 26400 104 26440
rect -396 26040 104 26080
rect -396 25620 -356 26040
rect 64 25620 104 26040
rect -396 25580 104 25620
rect -396 25220 104 25260
rect -396 24800 -356 25220
rect 64 24800 104 25220
rect -396 24760 104 24800
rect -396 24400 104 24440
rect -396 23980 -356 24400
rect 64 23980 104 24400
rect -396 23940 104 23980
rect -396 23580 104 23620
rect -396 23160 -356 23580
rect 64 23160 104 23580
rect -396 23120 104 23160
rect -396 22760 104 22800
rect -396 22340 -356 22760
rect 64 22340 104 22760
rect -396 22300 104 22340
rect -396 21940 104 21980
rect -396 21520 -356 21940
rect 64 21520 104 21940
rect -396 21480 104 21520
rect -396 21120 104 21160
rect -396 20700 -356 21120
rect 64 20700 104 21120
rect -396 20660 104 20700
rect -396 20300 104 20340
rect -396 19880 -356 20300
rect 64 19880 104 20300
rect -396 19840 104 19880
rect -396 19480 104 19520
rect -396 19060 -356 19480
rect 64 19060 104 19480
rect -396 19020 104 19060
rect -396 18660 104 18700
rect -396 18240 -356 18660
rect 64 18240 104 18660
rect -396 18200 104 18240
rect -396 17840 104 17880
rect -396 17420 -356 17840
rect 64 17420 104 17840
rect -396 17380 104 17420
rect -396 17020 104 17060
rect -396 16600 -356 17020
rect 64 16600 104 17020
rect -396 16560 104 16600
rect -396 16200 104 16240
rect -396 15780 -356 16200
rect 64 15780 104 16200
rect -396 15740 104 15780
rect -396 15380 104 15420
rect -396 14960 -356 15380
rect 64 14960 104 15380
rect -396 14920 104 14960
rect -396 14560 104 14600
rect -396 14140 -356 14560
rect 64 14140 104 14560
rect -396 14100 104 14140
rect -396 13740 104 13780
rect -396 13320 -356 13740
rect 64 13320 104 13740
rect -396 13280 104 13320
rect -396 12920 104 12960
rect -396 12500 -356 12920
rect 64 12500 104 12920
rect -396 12460 104 12500
rect -396 12100 104 12140
rect -396 11680 -356 12100
rect 64 11680 104 12100
rect -396 11640 104 11680
rect -396 11280 104 11320
rect -396 10860 -356 11280
rect 64 10860 104 11280
rect -396 10820 104 10860
rect -396 10460 104 10500
rect -396 10040 -356 10460
rect 64 10040 104 10460
rect -396 10000 104 10040
rect -396 9640 104 9680
rect -396 9220 -356 9640
rect 64 9220 104 9640
rect -396 9180 104 9220
rect -396 8820 104 8860
rect -396 8400 -356 8820
rect 64 8400 104 8820
rect -396 8360 104 8400
rect -396 8000 104 8040
rect -396 7580 -356 8000
rect 64 7580 104 8000
rect -396 7540 104 7580
rect -396 7180 104 7220
rect -396 6760 -356 7180
rect 64 6760 104 7180
rect -396 6720 104 6760
rect -396 6360 104 6400
rect -396 5940 -356 6360
rect 64 5940 104 6360
rect -396 5900 104 5940
rect -396 5540 104 5580
rect -396 5120 -356 5540
rect 64 5120 104 5540
rect -396 5080 104 5120
rect -396 4720 104 4760
rect -396 4300 -356 4720
rect 64 4300 104 4720
rect -396 4260 104 4300
rect -396 3900 104 3940
rect -396 3480 -356 3900
rect 64 3480 104 3900
rect -396 3440 104 3480
rect -396 3080 104 3120
rect -396 2660 -356 3080
rect 64 2660 104 3080
rect -396 2620 104 2660
rect -396 2260 104 2300
rect -396 1840 -356 2260
rect 64 1840 104 2260
rect -396 1800 104 1840
rect -396 1440 104 1480
rect -396 1020 -356 1440
rect 64 1020 104 1440
rect -396 980 104 1020
rect -396 620 104 660
rect -396 200 -356 620
rect 64 200 104 620
rect -396 160 104 200
rect -396 -200 104 -160
rect -396 -620 -356 -200
rect 64 -620 104 -200
rect -396 -660 104 -620
rect -396 -1020 104 -980
rect -396 -1440 -356 -1020
rect 64 -1440 104 -1020
rect -396 -1480 104 -1440
rect -396 -1840 104 -1800
rect -396 -2260 -356 -1840
rect 64 -2260 104 -1840
rect -396 -2300 104 -2260
rect -396 -2660 104 -2620
rect -396 -3080 -356 -2660
rect 64 -3080 104 -2660
rect -396 -3120 104 -3080
rect -396 -3480 104 -3440
rect -396 -3900 -356 -3480
rect 64 -3900 104 -3480
rect -396 -3940 104 -3900
rect -396 -4300 104 -4260
rect -396 -4720 -356 -4300
rect 64 -4720 104 -4300
rect -396 -4760 104 -4720
rect -396 -5120 104 -5080
rect -396 -5540 -356 -5120
rect 64 -5540 104 -5120
rect -396 -5580 104 -5540
rect -396 -5940 104 -5900
rect -396 -6360 -356 -5940
rect 64 -6360 104 -5940
rect -396 -6400 104 -6360
rect -396 -6760 104 -6720
rect -396 -7180 -356 -6760
rect 64 -7180 104 -6760
rect -396 -7220 104 -7180
rect -396 -7580 104 -7540
rect -396 -8000 -356 -7580
rect 64 -8000 104 -7580
rect -396 -8040 104 -8000
rect -396 -8400 104 -8360
rect -396 -8820 -356 -8400
rect 64 -8820 104 -8400
rect -396 -8860 104 -8820
rect -396 -9220 104 -9180
rect -396 -9640 -356 -9220
rect 64 -9640 104 -9220
rect -396 -9680 104 -9640
rect -396 -10040 104 -10000
rect -396 -10460 -356 -10040
rect 64 -10460 104 -10040
rect -396 -10500 104 -10460
rect -396 -10860 104 -10820
rect -396 -11280 -356 -10860
rect 64 -11280 104 -10860
rect -396 -11320 104 -11280
rect -396 -11680 104 -11640
rect -396 -12100 -356 -11680
rect 64 -12100 104 -11680
rect -396 -12140 104 -12100
rect -396 -12500 104 -12460
rect -396 -12920 -356 -12500
rect 64 -12920 104 -12500
rect -396 -12960 104 -12920
rect -396 -13320 104 -13280
rect -396 -13740 -356 -13320
rect 64 -13740 104 -13320
rect -396 -13780 104 -13740
rect -396 -14140 104 -14100
rect -396 -14560 -356 -14140
rect 64 -14560 104 -14140
rect -396 -14600 104 -14560
rect -396 -14960 104 -14920
rect -396 -15380 -356 -14960
rect 64 -15380 104 -14960
rect -396 -15420 104 -15380
rect -396 -15780 104 -15740
rect -396 -16200 -356 -15780
rect 64 -16200 104 -15780
rect -396 -16240 104 -16200
rect -396 -16600 104 -16560
rect -396 -17020 -356 -16600
rect 64 -17020 104 -16600
rect -396 -17060 104 -17020
rect -396 -17420 104 -17380
rect -396 -17840 -356 -17420
rect 64 -17840 104 -17420
rect -396 -17880 104 -17840
rect -396 -18240 104 -18200
rect -396 -18660 -356 -18240
rect 64 -18660 104 -18240
rect -396 -18700 104 -18660
rect -396 -19060 104 -19020
rect -396 -19480 -356 -19060
rect 64 -19480 104 -19060
rect -396 -19520 104 -19480
rect -396 -19880 104 -19840
rect -396 -20300 -356 -19880
rect 64 -20300 104 -19880
rect -396 -20340 104 -20300
rect -396 -20700 104 -20660
rect -396 -21120 -356 -20700
rect 64 -21120 104 -20700
rect -396 -21160 104 -21120
rect -396 -21520 104 -21480
rect -396 -21940 -356 -21520
rect 64 -21940 104 -21520
rect -396 -21980 104 -21940
rect -396 -22340 104 -22300
rect -396 -22760 -356 -22340
rect 64 -22760 104 -22340
rect -396 -22800 104 -22760
rect -396 -23160 104 -23120
rect -396 -23580 -356 -23160
rect 64 -23580 104 -23160
rect -396 -23620 104 -23580
rect -396 -23980 104 -23940
rect -396 -24400 -356 -23980
rect 64 -24400 104 -23980
rect -396 -24440 104 -24400
rect -396 -24800 104 -24760
rect -396 -25220 -356 -24800
rect 64 -25220 104 -24800
rect -396 -25260 104 -25220
rect -396 -25620 104 -25580
rect -396 -26040 -356 -25620
rect 64 -26040 104 -25620
rect -396 -26080 104 -26040
rect -396 -26440 104 -26400
rect -396 -26860 -356 -26440
rect 64 -26860 104 -26440
rect -396 -26900 104 -26860
rect -396 -27260 104 -27220
rect -396 -27680 -356 -27260
rect 64 -27680 104 -27260
rect -396 -27720 104 -27680
rect -396 -28080 104 -28040
rect -396 -28500 -356 -28080
rect 64 -28500 104 -28080
rect -396 -28540 104 -28500
rect -396 -28900 104 -28860
rect -396 -29320 -356 -28900
rect 64 -29320 104 -28900
rect -396 -29360 104 -29320
rect -396 -29720 104 -29680
rect -396 -30140 -356 -29720
rect 64 -30140 104 -29720
rect -396 -30180 104 -30140
rect -396 -30540 104 -30500
rect -396 -30960 -356 -30540
rect 64 -30960 104 -30540
rect -396 -31000 104 -30960
rect -396 -31360 104 -31320
rect -396 -31780 -356 -31360
rect 64 -31780 104 -31360
rect -396 -31820 104 -31780
rect -396 -32180 104 -32140
rect -396 -32600 -356 -32180
rect 64 -32600 104 -32180
rect -396 -32640 104 -32600
rect -396 -33000 104 -32960
rect -396 -33420 -356 -33000
rect 64 -33420 104 -33000
rect -396 -33460 104 -33420
rect -396 -33820 104 -33780
rect -396 -34240 -356 -33820
rect 64 -34240 104 -33820
rect -396 -34280 104 -34240
rect -396 -34640 104 -34600
rect -396 -35060 -356 -34640
rect 64 -35060 104 -34640
rect -396 -35100 104 -35060
rect -396 -35460 104 -35420
rect -396 -35880 -356 -35460
rect 64 -35880 104 -35460
rect -396 -35920 104 -35880
rect -396 -36280 104 -36240
rect -396 -36700 -356 -36280
rect 64 -36700 104 -36280
rect -396 -36740 104 -36700
rect -396 -37100 104 -37060
rect -396 -37520 -356 -37100
rect 64 -37520 104 -37100
rect -396 -37560 104 -37520
rect -396 -37920 104 -37880
rect -396 -38340 -356 -37920
rect 64 -38340 104 -37920
rect -396 -38380 104 -38340
rect -396 -38740 104 -38700
rect -396 -39160 -356 -38740
rect 64 -39160 104 -38740
rect -396 -39200 104 -39160
rect -396 -39560 104 -39520
rect -396 -39980 -356 -39560
rect 64 -39980 104 -39560
rect -396 -40020 104 -39980
rect -396 -40380 104 -40340
rect -396 -40800 -356 -40380
rect 64 -40800 104 -40380
rect -396 -40840 104 -40800
<< mimcapcontact >>
rect -356 40380 64 40800
rect -356 39560 64 39980
rect -356 38740 64 39160
rect -356 37920 64 38340
rect -356 37100 64 37520
rect -356 36280 64 36700
rect -356 35460 64 35880
rect -356 34640 64 35060
rect -356 33820 64 34240
rect -356 33000 64 33420
rect -356 32180 64 32600
rect -356 31360 64 31780
rect -356 30540 64 30960
rect -356 29720 64 30140
rect -356 28900 64 29320
rect -356 28080 64 28500
rect -356 27260 64 27680
rect -356 26440 64 26860
rect -356 25620 64 26040
rect -356 24800 64 25220
rect -356 23980 64 24400
rect -356 23160 64 23580
rect -356 22340 64 22760
rect -356 21520 64 21940
rect -356 20700 64 21120
rect -356 19880 64 20300
rect -356 19060 64 19480
rect -356 18240 64 18660
rect -356 17420 64 17840
rect -356 16600 64 17020
rect -356 15780 64 16200
rect -356 14960 64 15380
rect -356 14140 64 14560
rect -356 13320 64 13740
rect -356 12500 64 12920
rect -356 11680 64 12100
rect -356 10860 64 11280
rect -356 10040 64 10460
rect -356 9220 64 9640
rect -356 8400 64 8820
rect -356 7580 64 8000
rect -356 6760 64 7180
rect -356 5940 64 6360
rect -356 5120 64 5540
rect -356 4300 64 4720
rect -356 3480 64 3900
rect -356 2660 64 3080
rect -356 1840 64 2260
rect -356 1020 64 1440
rect -356 200 64 620
rect -356 -620 64 -200
rect -356 -1440 64 -1020
rect -356 -2260 64 -1840
rect -356 -3080 64 -2660
rect -356 -3900 64 -3480
rect -356 -4720 64 -4300
rect -356 -5540 64 -5120
rect -356 -6360 64 -5940
rect -356 -7180 64 -6760
rect -356 -8000 64 -7580
rect -356 -8820 64 -8400
rect -356 -9640 64 -9220
rect -356 -10460 64 -10040
rect -356 -11280 64 -10860
rect -356 -12100 64 -11680
rect -356 -12920 64 -12500
rect -356 -13740 64 -13320
rect -356 -14560 64 -14140
rect -356 -15380 64 -14960
rect -356 -16200 64 -15780
rect -356 -17020 64 -16600
rect -356 -17840 64 -17420
rect -356 -18660 64 -18240
rect -356 -19480 64 -19060
rect -356 -20300 64 -19880
rect -356 -21120 64 -20700
rect -356 -21940 64 -21520
rect -356 -22760 64 -22340
rect -356 -23580 64 -23160
rect -356 -24400 64 -23980
rect -356 -25220 64 -24800
rect -356 -26040 64 -25620
rect -356 -26860 64 -26440
rect -356 -27680 64 -27260
rect -356 -28500 64 -28080
rect -356 -29320 64 -28900
rect -356 -30140 64 -29720
rect -356 -30960 64 -30540
rect -356 -31780 64 -31360
rect -356 -32600 64 -32180
rect -356 -33420 64 -33000
rect -356 -34240 64 -33820
rect -356 -35060 64 -34640
rect -356 -35880 64 -35460
rect -356 -36700 64 -36280
rect -356 -37520 64 -37100
rect -356 -38340 64 -37920
rect -356 -39160 64 -38740
rect -356 -39980 64 -39560
rect -356 -40800 64 -40380
<< metal4 >>
rect -198 40801 -94 41000
rect 332 40852 436 41000
rect -357 40800 65 40801
rect -357 40380 -356 40800
rect 64 40380 65 40800
rect -357 40379 65 40380
rect -198 39981 -94 40379
rect 332 40328 352 40852
rect 416 40328 436 40852
rect 332 40032 436 40328
rect -357 39980 65 39981
rect -357 39560 -356 39980
rect 64 39560 65 39980
rect -357 39559 65 39560
rect -198 39161 -94 39559
rect 332 39508 352 40032
rect 416 39508 436 40032
rect 332 39212 436 39508
rect -357 39160 65 39161
rect -357 38740 -356 39160
rect 64 38740 65 39160
rect -357 38739 65 38740
rect -198 38341 -94 38739
rect 332 38688 352 39212
rect 416 38688 436 39212
rect 332 38392 436 38688
rect -357 38340 65 38341
rect -357 37920 -356 38340
rect 64 37920 65 38340
rect -357 37919 65 37920
rect -198 37521 -94 37919
rect 332 37868 352 38392
rect 416 37868 436 38392
rect 332 37572 436 37868
rect -357 37520 65 37521
rect -357 37100 -356 37520
rect 64 37100 65 37520
rect -357 37099 65 37100
rect -198 36701 -94 37099
rect 332 37048 352 37572
rect 416 37048 436 37572
rect 332 36752 436 37048
rect -357 36700 65 36701
rect -357 36280 -356 36700
rect 64 36280 65 36700
rect -357 36279 65 36280
rect -198 35881 -94 36279
rect 332 36228 352 36752
rect 416 36228 436 36752
rect 332 35932 436 36228
rect -357 35880 65 35881
rect -357 35460 -356 35880
rect 64 35460 65 35880
rect -357 35459 65 35460
rect -198 35061 -94 35459
rect 332 35408 352 35932
rect 416 35408 436 35932
rect 332 35112 436 35408
rect -357 35060 65 35061
rect -357 34640 -356 35060
rect 64 34640 65 35060
rect -357 34639 65 34640
rect -198 34241 -94 34639
rect 332 34588 352 35112
rect 416 34588 436 35112
rect 332 34292 436 34588
rect -357 34240 65 34241
rect -357 33820 -356 34240
rect 64 33820 65 34240
rect -357 33819 65 33820
rect -198 33421 -94 33819
rect 332 33768 352 34292
rect 416 33768 436 34292
rect 332 33472 436 33768
rect -357 33420 65 33421
rect -357 33000 -356 33420
rect 64 33000 65 33420
rect -357 32999 65 33000
rect -198 32601 -94 32999
rect 332 32948 352 33472
rect 416 32948 436 33472
rect 332 32652 436 32948
rect -357 32600 65 32601
rect -357 32180 -356 32600
rect 64 32180 65 32600
rect -357 32179 65 32180
rect -198 31781 -94 32179
rect 332 32128 352 32652
rect 416 32128 436 32652
rect 332 31832 436 32128
rect -357 31780 65 31781
rect -357 31360 -356 31780
rect 64 31360 65 31780
rect -357 31359 65 31360
rect -198 30961 -94 31359
rect 332 31308 352 31832
rect 416 31308 436 31832
rect 332 31012 436 31308
rect -357 30960 65 30961
rect -357 30540 -356 30960
rect 64 30540 65 30960
rect -357 30539 65 30540
rect -198 30141 -94 30539
rect 332 30488 352 31012
rect 416 30488 436 31012
rect 332 30192 436 30488
rect -357 30140 65 30141
rect -357 29720 -356 30140
rect 64 29720 65 30140
rect -357 29719 65 29720
rect -198 29321 -94 29719
rect 332 29668 352 30192
rect 416 29668 436 30192
rect 332 29372 436 29668
rect -357 29320 65 29321
rect -357 28900 -356 29320
rect 64 28900 65 29320
rect -357 28899 65 28900
rect -198 28501 -94 28899
rect 332 28848 352 29372
rect 416 28848 436 29372
rect 332 28552 436 28848
rect -357 28500 65 28501
rect -357 28080 -356 28500
rect 64 28080 65 28500
rect -357 28079 65 28080
rect -198 27681 -94 28079
rect 332 28028 352 28552
rect 416 28028 436 28552
rect 332 27732 436 28028
rect -357 27680 65 27681
rect -357 27260 -356 27680
rect 64 27260 65 27680
rect -357 27259 65 27260
rect -198 26861 -94 27259
rect 332 27208 352 27732
rect 416 27208 436 27732
rect 332 26912 436 27208
rect -357 26860 65 26861
rect -357 26440 -356 26860
rect 64 26440 65 26860
rect -357 26439 65 26440
rect -198 26041 -94 26439
rect 332 26388 352 26912
rect 416 26388 436 26912
rect 332 26092 436 26388
rect -357 26040 65 26041
rect -357 25620 -356 26040
rect 64 25620 65 26040
rect -357 25619 65 25620
rect -198 25221 -94 25619
rect 332 25568 352 26092
rect 416 25568 436 26092
rect 332 25272 436 25568
rect -357 25220 65 25221
rect -357 24800 -356 25220
rect 64 24800 65 25220
rect -357 24799 65 24800
rect -198 24401 -94 24799
rect 332 24748 352 25272
rect 416 24748 436 25272
rect 332 24452 436 24748
rect -357 24400 65 24401
rect -357 23980 -356 24400
rect 64 23980 65 24400
rect -357 23979 65 23980
rect -198 23581 -94 23979
rect 332 23928 352 24452
rect 416 23928 436 24452
rect 332 23632 436 23928
rect -357 23580 65 23581
rect -357 23160 -356 23580
rect 64 23160 65 23580
rect -357 23159 65 23160
rect -198 22761 -94 23159
rect 332 23108 352 23632
rect 416 23108 436 23632
rect 332 22812 436 23108
rect -357 22760 65 22761
rect -357 22340 -356 22760
rect 64 22340 65 22760
rect -357 22339 65 22340
rect -198 21941 -94 22339
rect 332 22288 352 22812
rect 416 22288 436 22812
rect 332 21992 436 22288
rect -357 21940 65 21941
rect -357 21520 -356 21940
rect 64 21520 65 21940
rect -357 21519 65 21520
rect -198 21121 -94 21519
rect 332 21468 352 21992
rect 416 21468 436 21992
rect 332 21172 436 21468
rect -357 21120 65 21121
rect -357 20700 -356 21120
rect 64 20700 65 21120
rect -357 20699 65 20700
rect -198 20301 -94 20699
rect 332 20648 352 21172
rect 416 20648 436 21172
rect 332 20352 436 20648
rect -357 20300 65 20301
rect -357 19880 -356 20300
rect 64 19880 65 20300
rect -357 19879 65 19880
rect -198 19481 -94 19879
rect 332 19828 352 20352
rect 416 19828 436 20352
rect 332 19532 436 19828
rect -357 19480 65 19481
rect -357 19060 -356 19480
rect 64 19060 65 19480
rect -357 19059 65 19060
rect -198 18661 -94 19059
rect 332 19008 352 19532
rect 416 19008 436 19532
rect 332 18712 436 19008
rect -357 18660 65 18661
rect -357 18240 -356 18660
rect 64 18240 65 18660
rect -357 18239 65 18240
rect -198 17841 -94 18239
rect 332 18188 352 18712
rect 416 18188 436 18712
rect 332 17892 436 18188
rect -357 17840 65 17841
rect -357 17420 -356 17840
rect 64 17420 65 17840
rect -357 17419 65 17420
rect -198 17021 -94 17419
rect 332 17368 352 17892
rect 416 17368 436 17892
rect 332 17072 436 17368
rect -357 17020 65 17021
rect -357 16600 -356 17020
rect 64 16600 65 17020
rect -357 16599 65 16600
rect -198 16201 -94 16599
rect 332 16548 352 17072
rect 416 16548 436 17072
rect 332 16252 436 16548
rect -357 16200 65 16201
rect -357 15780 -356 16200
rect 64 15780 65 16200
rect -357 15779 65 15780
rect -198 15381 -94 15779
rect 332 15728 352 16252
rect 416 15728 436 16252
rect 332 15432 436 15728
rect -357 15380 65 15381
rect -357 14960 -356 15380
rect 64 14960 65 15380
rect -357 14959 65 14960
rect -198 14561 -94 14959
rect 332 14908 352 15432
rect 416 14908 436 15432
rect 332 14612 436 14908
rect -357 14560 65 14561
rect -357 14140 -356 14560
rect 64 14140 65 14560
rect -357 14139 65 14140
rect -198 13741 -94 14139
rect 332 14088 352 14612
rect 416 14088 436 14612
rect 332 13792 436 14088
rect -357 13740 65 13741
rect -357 13320 -356 13740
rect 64 13320 65 13740
rect -357 13319 65 13320
rect -198 12921 -94 13319
rect 332 13268 352 13792
rect 416 13268 436 13792
rect 332 12972 436 13268
rect -357 12920 65 12921
rect -357 12500 -356 12920
rect 64 12500 65 12920
rect -357 12499 65 12500
rect -198 12101 -94 12499
rect 332 12448 352 12972
rect 416 12448 436 12972
rect 332 12152 436 12448
rect -357 12100 65 12101
rect -357 11680 -356 12100
rect 64 11680 65 12100
rect -357 11679 65 11680
rect -198 11281 -94 11679
rect 332 11628 352 12152
rect 416 11628 436 12152
rect 332 11332 436 11628
rect -357 11280 65 11281
rect -357 10860 -356 11280
rect 64 10860 65 11280
rect -357 10859 65 10860
rect -198 10461 -94 10859
rect 332 10808 352 11332
rect 416 10808 436 11332
rect 332 10512 436 10808
rect -357 10460 65 10461
rect -357 10040 -356 10460
rect 64 10040 65 10460
rect -357 10039 65 10040
rect -198 9641 -94 10039
rect 332 9988 352 10512
rect 416 9988 436 10512
rect 332 9692 436 9988
rect -357 9640 65 9641
rect -357 9220 -356 9640
rect 64 9220 65 9640
rect -357 9219 65 9220
rect -198 8821 -94 9219
rect 332 9168 352 9692
rect 416 9168 436 9692
rect 332 8872 436 9168
rect -357 8820 65 8821
rect -357 8400 -356 8820
rect 64 8400 65 8820
rect -357 8399 65 8400
rect -198 8001 -94 8399
rect 332 8348 352 8872
rect 416 8348 436 8872
rect 332 8052 436 8348
rect -357 8000 65 8001
rect -357 7580 -356 8000
rect 64 7580 65 8000
rect -357 7579 65 7580
rect -198 7181 -94 7579
rect 332 7528 352 8052
rect 416 7528 436 8052
rect 332 7232 436 7528
rect -357 7180 65 7181
rect -357 6760 -356 7180
rect 64 6760 65 7180
rect -357 6759 65 6760
rect -198 6361 -94 6759
rect 332 6708 352 7232
rect 416 6708 436 7232
rect 332 6412 436 6708
rect -357 6360 65 6361
rect -357 5940 -356 6360
rect 64 5940 65 6360
rect -357 5939 65 5940
rect -198 5541 -94 5939
rect 332 5888 352 6412
rect 416 5888 436 6412
rect 332 5592 436 5888
rect -357 5540 65 5541
rect -357 5120 -356 5540
rect 64 5120 65 5540
rect -357 5119 65 5120
rect -198 4721 -94 5119
rect 332 5068 352 5592
rect 416 5068 436 5592
rect 332 4772 436 5068
rect -357 4720 65 4721
rect -357 4300 -356 4720
rect 64 4300 65 4720
rect -357 4299 65 4300
rect -198 3901 -94 4299
rect 332 4248 352 4772
rect 416 4248 436 4772
rect 332 3952 436 4248
rect -357 3900 65 3901
rect -357 3480 -356 3900
rect 64 3480 65 3900
rect -357 3479 65 3480
rect -198 3081 -94 3479
rect 332 3428 352 3952
rect 416 3428 436 3952
rect 332 3132 436 3428
rect -357 3080 65 3081
rect -357 2660 -356 3080
rect 64 2660 65 3080
rect -357 2659 65 2660
rect -198 2261 -94 2659
rect 332 2608 352 3132
rect 416 2608 436 3132
rect 332 2312 436 2608
rect -357 2260 65 2261
rect -357 1840 -356 2260
rect 64 1840 65 2260
rect -357 1839 65 1840
rect -198 1441 -94 1839
rect 332 1788 352 2312
rect 416 1788 436 2312
rect 332 1492 436 1788
rect -357 1440 65 1441
rect -357 1020 -356 1440
rect 64 1020 65 1440
rect -357 1019 65 1020
rect -198 621 -94 1019
rect 332 968 352 1492
rect 416 968 436 1492
rect 332 672 436 968
rect -357 620 65 621
rect -357 200 -356 620
rect 64 200 65 620
rect -357 199 65 200
rect -198 -199 -94 199
rect 332 148 352 672
rect 416 148 436 672
rect 332 -148 436 148
rect -357 -200 65 -199
rect -357 -620 -356 -200
rect 64 -620 65 -200
rect -357 -621 65 -620
rect -198 -1019 -94 -621
rect 332 -672 352 -148
rect 416 -672 436 -148
rect 332 -968 436 -672
rect -357 -1020 65 -1019
rect -357 -1440 -356 -1020
rect 64 -1440 65 -1020
rect -357 -1441 65 -1440
rect -198 -1839 -94 -1441
rect 332 -1492 352 -968
rect 416 -1492 436 -968
rect 332 -1788 436 -1492
rect -357 -1840 65 -1839
rect -357 -2260 -356 -1840
rect 64 -2260 65 -1840
rect -357 -2261 65 -2260
rect -198 -2659 -94 -2261
rect 332 -2312 352 -1788
rect 416 -2312 436 -1788
rect 332 -2608 436 -2312
rect -357 -2660 65 -2659
rect -357 -3080 -356 -2660
rect 64 -3080 65 -2660
rect -357 -3081 65 -3080
rect -198 -3479 -94 -3081
rect 332 -3132 352 -2608
rect 416 -3132 436 -2608
rect 332 -3428 436 -3132
rect -357 -3480 65 -3479
rect -357 -3900 -356 -3480
rect 64 -3900 65 -3480
rect -357 -3901 65 -3900
rect -198 -4299 -94 -3901
rect 332 -3952 352 -3428
rect 416 -3952 436 -3428
rect 332 -4248 436 -3952
rect -357 -4300 65 -4299
rect -357 -4720 -356 -4300
rect 64 -4720 65 -4300
rect -357 -4721 65 -4720
rect -198 -5119 -94 -4721
rect 332 -4772 352 -4248
rect 416 -4772 436 -4248
rect 332 -5068 436 -4772
rect -357 -5120 65 -5119
rect -357 -5540 -356 -5120
rect 64 -5540 65 -5120
rect -357 -5541 65 -5540
rect -198 -5939 -94 -5541
rect 332 -5592 352 -5068
rect 416 -5592 436 -5068
rect 332 -5888 436 -5592
rect -357 -5940 65 -5939
rect -357 -6360 -356 -5940
rect 64 -6360 65 -5940
rect -357 -6361 65 -6360
rect -198 -6759 -94 -6361
rect 332 -6412 352 -5888
rect 416 -6412 436 -5888
rect 332 -6708 436 -6412
rect -357 -6760 65 -6759
rect -357 -7180 -356 -6760
rect 64 -7180 65 -6760
rect -357 -7181 65 -7180
rect -198 -7579 -94 -7181
rect 332 -7232 352 -6708
rect 416 -7232 436 -6708
rect 332 -7528 436 -7232
rect -357 -7580 65 -7579
rect -357 -8000 -356 -7580
rect 64 -8000 65 -7580
rect -357 -8001 65 -8000
rect -198 -8399 -94 -8001
rect 332 -8052 352 -7528
rect 416 -8052 436 -7528
rect 332 -8348 436 -8052
rect -357 -8400 65 -8399
rect -357 -8820 -356 -8400
rect 64 -8820 65 -8400
rect -357 -8821 65 -8820
rect -198 -9219 -94 -8821
rect 332 -8872 352 -8348
rect 416 -8872 436 -8348
rect 332 -9168 436 -8872
rect -357 -9220 65 -9219
rect -357 -9640 -356 -9220
rect 64 -9640 65 -9220
rect -357 -9641 65 -9640
rect -198 -10039 -94 -9641
rect 332 -9692 352 -9168
rect 416 -9692 436 -9168
rect 332 -9988 436 -9692
rect -357 -10040 65 -10039
rect -357 -10460 -356 -10040
rect 64 -10460 65 -10040
rect -357 -10461 65 -10460
rect -198 -10859 -94 -10461
rect 332 -10512 352 -9988
rect 416 -10512 436 -9988
rect 332 -10808 436 -10512
rect -357 -10860 65 -10859
rect -357 -11280 -356 -10860
rect 64 -11280 65 -10860
rect -357 -11281 65 -11280
rect -198 -11679 -94 -11281
rect 332 -11332 352 -10808
rect 416 -11332 436 -10808
rect 332 -11628 436 -11332
rect -357 -11680 65 -11679
rect -357 -12100 -356 -11680
rect 64 -12100 65 -11680
rect -357 -12101 65 -12100
rect -198 -12499 -94 -12101
rect 332 -12152 352 -11628
rect 416 -12152 436 -11628
rect 332 -12448 436 -12152
rect -357 -12500 65 -12499
rect -357 -12920 -356 -12500
rect 64 -12920 65 -12500
rect -357 -12921 65 -12920
rect -198 -13319 -94 -12921
rect 332 -12972 352 -12448
rect 416 -12972 436 -12448
rect 332 -13268 436 -12972
rect -357 -13320 65 -13319
rect -357 -13740 -356 -13320
rect 64 -13740 65 -13320
rect -357 -13741 65 -13740
rect -198 -14139 -94 -13741
rect 332 -13792 352 -13268
rect 416 -13792 436 -13268
rect 332 -14088 436 -13792
rect -357 -14140 65 -14139
rect -357 -14560 -356 -14140
rect 64 -14560 65 -14140
rect -357 -14561 65 -14560
rect -198 -14959 -94 -14561
rect 332 -14612 352 -14088
rect 416 -14612 436 -14088
rect 332 -14908 436 -14612
rect -357 -14960 65 -14959
rect -357 -15380 -356 -14960
rect 64 -15380 65 -14960
rect -357 -15381 65 -15380
rect -198 -15779 -94 -15381
rect 332 -15432 352 -14908
rect 416 -15432 436 -14908
rect 332 -15728 436 -15432
rect -357 -15780 65 -15779
rect -357 -16200 -356 -15780
rect 64 -16200 65 -15780
rect -357 -16201 65 -16200
rect -198 -16599 -94 -16201
rect 332 -16252 352 -15728
rect 416 -16252 436 -15728
rect 332 -16548 436 -16252
rect -357 -16600 65 -16599
rect -357 -17020 -356 -16600
rect 64 -17020 65 -16600
rect -357 -17021 65 -17020
rect -198 -17419 -94 -17021
rect 332 -17072 352 -16548
rect 416 -17072 436 -16548
rect 332 -17368 436 -17072
rect -357 -17420 65 -17419
rect -357 -17840 -356 -17420
rect 64 -17840 65 -17420
rect -357 -17841 65 -17840
rect -198 -18239 -94 -17841
rect 332 -17892 352 -17368
rect 416 -17892 436 -17368
rect 332 -18188 436 -17892
rect -357 -18240 65 -18239
rect -357 -18660 -356 -18240
rect 64 -18660 65 -18240
rect -357 -18661 65 -18660
rect -198 -19059 -94 -18661
rect 332 -18712 352 -18188
rect 416 -18712 436 -18188
rect 332 -19008 436 -18712
rect -357 -19060 65 -19059
rect -357 -19480 -356 -19060
rect 64 -19480 65 -19060
rect -357 -19481 65 -19480
rect -198 -19879 -94 -19481
rect 332 -19532 352 -19008
rect 416 -19532 436 -19008
rect 332 -19828 436 -19532
rect -357 -19880 65 -19879
rect -357 -20300 -356 -19880
rect 64 -20300 65 -19880
rect -357 -20301 65 -20300
rect -198 -20699 -94 -20301
rect 332 -20352 352 -19828
rect 416 -20352 436 -19828
rect 332 -20648 436 -20352
rect -357 -20700 65 -20699
rect -357 -21120 -356 -20700
rect 64 -21120 65 -20700
rect -357 -21121 65 -21120
rect -198 -21519 -94 -21121
rect 332 -21172 352 -20648
rect 416 -21172 436 -20648
rect 332 -21468 436 -21172
rect -357 -21520 65 -21519
rect -357 -21940 -356 -21520
rect 64 -21940 65 -21520
rect -357 -21941 65 -21940
rect -198 -22339 -94 -21941
rect 332 -21992 352 -21468
rect 416 -21992 436 -21468
rect 332 -22288 436 -21992
rect -357 -22340 65 -22339
rect -357 -22760 -356 -22340
rect 64 -22760 65 -22340
rect -357 -22761 65 -22760
rect -198 -23159 -94 -22761
rect 332 -22812 352 -22288
rect 416 -22812 436 -22288
rect 332 -23108 436 -22812
rect -357 -23160 65 -23159
rect -357 -23580 -356 -23160
rect 64 -23580 65 -23160
rect -357 -23581 65 -23580
rect -198 -23979 -94 -23581
rect 332 -23632 352 -23108
rect 416 -23632 436 -23108
rect 332 -23928 436 -23632
rect -357 -23980 65 -23979
rect -357 -24400 -356 -23980
rect 64 -24400 65 -23980
rect -357 -24401 65 -24400
rect -198 -24799 -94 -24401
rect 332 -24452 352 -23928
rect 416 -24452 436 -23928
rect 332 -24748 436 -24452
rect -357 -24800 65 -24799
rect -357 -25220 -356 -24800
rect 64 -25220 65 -24800
rect -357 -25221 65 -25220
rect -198 -25619 -94 -25221
rect 332 -25272 352 -24748
rect 416 -25272 436 -24748
rect 332 -25568 436 -25272
rect -357 -25620 65 -25619
rect -357 -26040 -356 -25620
rect 64 -26040 65 -25620
rect -357 -26041 65 -26040
rect -198 -26439 -94 -26041
rect 332 -26092 352 -25568
rect 416 -26092 436 -25568
rect 332 -26388 436 -26092
rect -357 -26440 65 -26439
rect -357 -26860 -356 -26440
rect 64 -26860 65 -26440
rect -357 -26861 65 -26860
rect -198 -27259 -94 -26861
rect 332 -26912 352 -26388
rect 416 -26912 436 -26388
rect 332 -27208 436 -26912
rect -357 -27260 65 -27259
rect -357 -27680 -356 -27260
rect 64 -27680 65 -27260
rect -357 -27681 65 -27680
rect -198 -28079 -94 -27681
rect 332 -27732 352 -27208
rect 416 -27732 436 -27208
rect 332 -28028 436 -27732
rect -357 -28080 65 -28079
rect -357 -28500 -356 -28080
rect 64 -28500 65 -28080
rect -357 -28501 65 -28500
rect -198 -28899 -94 -28501
rect 332 -28552 352 -28028
rect 416 -28552 436 -28028
rect 332 -28848 436 -28552
rect -357 -28900 65 -28899
rect -357 -29320 -356 -28900
rect 64 -29320 65 -28900
rect -357 -29321 65 -29320
rect -198 -29719 -94 -29321
rect 332 -29372 352 -28848
rect 416 -29372 436 -28848
rect 332 -29668 436 -29372
rect -357 -29720 65 -29719
rect -357 -30140 -356 -29720
rect 64 -30140 65 -29720
rect -357 -30141 65 -30140
rect -198 -30539 -94 -30141
rect 332 -30192 352 -29668
rect 416 -30192 436 -29668
rect 332 -30488 436 -30192
rect -357 -30540 65 -30539
rect -357 -30960 -356 -30540
rect 64 -30960 65 -30540
rect -357 -30961 65 -30960
rect -198 -31359 -94 -30961
rect 332 -31012 352 -30488
rect 416 -31012 436 -30488
rect 332 -31308 436 -31012
rect -357 -31360 65 -31359
rect -357 -31780 -356 -31360
rect 64 -31780 65 -31360
rect -357 -31781 65 -31780
rect -198 -32179 -94 -31781
rect 332 -31832 352 -31308
rect 416 -31832 436 -31308
rect 332 -32128 436 -31832
rect -357 -32180 65 -32179
rect -357 -32600 -356 -32180
rect 64 -32600 65 -32180
rect -357 -32601 65 -32600
rect -198 -32999 -94 -32601
rect 332 -32652 352 -32128
rect 416 -32652 436 -32128
rect 332 -32948 436 -32652
rect -357 -33000 65 -32999
rect -357 -33420 -356 -33000
rect 64 -33420 65 -33000
rect -357 -33421 65 -33420
rect -198 -33819 -94 -33421
rect 332 -33472 352 -32948
rect 416 -33472 436 -32948
rect 332 -33768 436 -33472
rect -357 -33820 65 -33819
rect -357 -34240 -356 -33820
rect 64 -34240 65 -33820
rect -357 -34241 65 -34240
rect -198 -34639 -94 -34241
rect 332 -34292 352 -33768
rect 416 -34292 436 -33768
rect 332 -34588 436 -34292
rect -357 -34640 65 -34639
rect -357 -35060 -356 -34640
rect 64 -35060 65 -34640
rect -357 -35061 65 -35060
rect -198 -35459 -94 -35061
rect 332 -35112 352 -34588
rect 416 -35112 436 -34588
rect 332 -35408 436 -35112
rect -357 -35460 65 -35459
rect -357 -35880 -356 -35460
rect 64 -35880 65 -35460
rect -357 -35881 65 -35880
rect -198 -36279 -94 -35881
rect 332 -35932 352 -35408
rect 416 -35932 436 -35408
rect 332 -36228 436 -35932
rect -357 -36280 65 -36279
rect -357 -36700 -356 -36280
rect 64 -36700 65 -36280
rect -357 -36701 65 -36700
rect -198 -37099 -94 -36701
rect 332 -36752 352 -36228
rect 416 -36752 436 -36228
rect 332 -37048 436 -36752
rect -357 -37100 65 -37099
rect -357 -37520 -356 -37100
rect 64 -37520 65 -37100
rect -357 -37521 65 -37520
rect -198 -37919 -94 -37521
rect 332 -37572 352 -37048
rect 416 -37572 436 -37048
rect 332 -37868 436 -37572
rect -357 -37920 65 -37919
rect -357 -38340 -356 -37920
rect 64 -38340 65 -37920
rect -357 -38341 65 -38340
rect -198 -38739 -94 -38341
rect 332 -38392 352 -37868
rect 416 -38392 436 -37868
rect 332 -38688 436 -38392
rect -357 -38740 65 -38739
rect -357 -39160 -356 -38740
rect 64 -39160 65 -38740
rect -357 -39161 65 -39160
rect -198 -39559 -94 -39161
rect 332 -39212 352 -38688
rect 416 -39212 436 -38688
rect 332 -39508 436 -39212
rect -357 -39560 65 -39559
rect -357 -39980 -356 -39560
rect 64 -39980 65 -39560
rect -357 -39981 65 -39980
rect -198 -40379 -94 -39981
rect 332 -40032 352 -39508
rect 416 -40032 436 -39508
rect 332 -40328 436 -40032
rect -357 -40380 65 -40379
rect -357 -40800 -356 -40380
rect 64 -40800 65 -40380
rect -357 -40801 65 -40800
rect -198 -41000 -94 -40801
rect 332 -40852 352 -40328
rect 416 -40852 436 -40328
rect 332 -41000 436 -40852
<< properties >>
string FIXED_BBOX -436 40300 144 40880
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.5 l 2.5 val 14.4 carea 2.00 cperi 0.19 nx 1 ny 100 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
