magic
tech sky130A
timestamp 1725609876
<< metal1 >>
rect 100 12710 2395 12715
rect 100 12620 105 12710
rect 295 12620 2395 12710
rect 100 12615 2395 12620
rect 400 12520 2410 12525
rect 400 12430 405 12520
rect 595 12430 2410 12520
rect 400 12425 2410 12430
rect 3650 625 3750 7040
rect 4220 950 4320 7045
rect 4220 945 13340 950
rect 4220 855 13255 945
rect 13335 855 13340 945
rect 4220 850 13340 855
rect 3650 620 15270 625
rect 3650 530 15185 620
rect 15265 530 15270 620
rect 3650 525 15270 530
<< via1 >>
rect 4930 16315 5025 16405
rect 5420 16315 5510 16405
rect 8480 16315 8570 16405
rect 8970 16315 9060 16405
rect 105 12620 295 12710
rect 405 12430 595 12520
rect 4930 8565 5020 8655
rect 5420 8565 5510 8655
rect 8480 8565 8570 8655
rect 8970 8565 9060 8655
rect 13255 855 13335 945
rect 15185 530 15265 620
<< metal2 >>
rect 4925 16405 5030 16410
rect 4925 16315 4930 16405
rect 5025 16315 5030 16405
rect 4925 16310 5030 16315
rect 5415 16405 5515 16410
rect 5415 16315 5420 16405
rect 5510 16315 5515 16405
rect 5415 16310 5515 16315
rect 8475 16405 8575 16410
rect 8475 16315 8480 16405
rect 8570 16315 8575 16405
rect 8475 16310 8575 16315
rect 8965 16405 9065 16410
rect 8965 16315 8970 16405
rect 9060 16315 9065 16405
rect 8965 16310 9065 16315
rect 100 12710 300 12715
rect 100 12620 105 12710
rect 295 12620 300 12710
rect 100 12615 300 12620
rect 400 12520 600 12525
rect 400 12430 405 12520
rect 595 12430 600 12520
rect 400 12425 600 12430
rect 4925 8655 5025 8660
rect 4925 8565 4930 8655
rect 5020 8565 5025 8655
rect 4925 8560 5025 8565
rect 5415 8655 5515 8660
rect 5415 8565 5420 8655
rect 5510 8565 5515 8655
rect 5415 8560 5515 8565
rect 8475 8655 8575 8660
rect 8475 8565 8480 8655
rect 8570 8565 8575 8655
rect 8475 8560 8575 8565
rect 8965 8655 9065 8660
rect 8965 8565 8970 8655
rect 9060 8565 9065 8655
rect 8965 8560 9065 8565
rect 13250 945 13340 950
rect 13250 855 13255 945
rect 13335 855 13340 945
rect 13250 850 13340 855
rect 15180 620 15270 625
rect 15180 530 15185 620
rect 15265 530 15270 620
rect 15180 525 15270 530
<< via2 >>
rect 4930 16315 5025 16405
rect 5420 16315 5510 16405
rect 8480 16315 8570 16405
rect 8970 16315 9060 16405
rect 105 12620 295 12710
rect 405 12430 595 12520
rect 4930 8565 5020 8655
rect 5420 8565 5510 8655
rect 8480 8565 8570 8655
rect 8970 8565 9060 8655
rect 13255 855 13335 945
rect 15185 530 15265 620
<< metal3 >>
rect 4925 16405 5030 16410
rect 4925 16315 4930 16405
rect 5025 16315 5030 16405
rect 4925 16310 5030 16315
rect 5415 16405 5515 16410
rect 5415 16315 5420 16405
rect 5510 16315 5515 16405
rect 5415 16310 5515 16315
rect 8475 16405 8575 16410
rect 8475 16315 8480 16405
rect 8570 16315 8575 16405
rect 8475 16310 8575 16315
rect 8965 16405 9065 16410
rect 8965 16315 8970 16405
rect 9060 16315 9065 16405
rect 8965 16310 9065 16315
rect 100 12710 300 12715
rect 100 12620 105 12710
rect 295 12620 300 12710
rect 100 12615 300 12620
rect 400 12520 600 12525
rect 400 12430 405 12520
rect 595 12430 600 12520
rect 400 12425 600 12430
rect 4925 8655 5025 8660
rect 4925 8565 4930 8655
rect 5020 8565 5025 8655
rect 4925 8560 5025 8565
rect 5415 8655 5515 8660
rect 5415 8565 5420 8655
rect 5510 8565 5515 8655
rect 5415 8560 5515 8565
rect 8475 8655 8575 8660
rect 8475 8565 8480 8655
rect 8570 8565 8575 8655
rect 8475 8560 8575 8565
rect 8965 8655 9065 8660
rect 8965 8565 8970 8655
rect 9060 8565 9065 8655
rect 8965 8560 9065 8565
rect 13250 945 13340 950
rect 13250 855 13255 945
rect 13335 855 13340 945
rect 13250 850 13340 855
rect 15180 620 15270 625
rect 15180 530 15185 620
rect 15265 530 15270 620
rect 15180 525 15270 530
<< via3 >>
rect 4930 16315 5025 16405
rect 5420 16315 5510 16405
rect 8480 16315 8570 16405
rect 8970 16315 9060 16405
rect 105 12620 295 12710
rect 405 12430 595 12520
rect 4930 8565 5020 8655
rect 5420 8565 5510 8655
rect 8480 8565 8570 8655
rect 8970 8565 9060 8655
rect 13255 855 13335 945
rect 15185 530 15265 620
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 3067 22446 7237 22476
rect 3067 22076 3097 22446
rect 100 12710 300 22076
rect 100 12620 105 12710
rect 295 12620 300 12710
rect 100 500 300 12620
rect 400 22046 3097 22076
rect 400 12520 600 22046
rect 7483 17325 7513 22576
rect 4985 17295 7513 17325
rect 4985 16410 5015 17295
rect 7759 17125 7789 22576
rect 5465 17095 7789 17125
rect 8035 17145 8065 22576
rect 8311 17375 8341 22576
rect 8587 17680 8617 22576
rect 8863 17960 8893 22576
rect 9139 18210 9169 22576
rect 9415 18455 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 9415 18425 12225 18455
rect 9139 18180 11895 18210
rect 8863 17930 11635 17960
rect 8587 17650 11415 17680
rect 8311 17345 9015 17375
rect 8035 17115 8530 17145
rect 5465 16410 5495 17095
rect 8500 16410 8530 17115
rect 8985 16410 9015 17345
rect 4925 16405 5030 16410
rect 4925 16315 4930 16405
rect 5025 16315 5030 16405
rect 4925 16310 5030 16315
rect 5415 16405 5515 16410
rect 5415 16315 5420 16405
rect 5510 16315 5515 16405
rect 5415 16310 5515 16315
rect 8475 16405 8575 16410
rect 8475 16315 8480 16405
rect 8570 16315 8575 16405
rect 8475 16310 8575 16315
rect 8965 16405 9065 16410
rect 8965 16315 8970 16405
rect 9060 16315 9065 16405
rect 8965 16310 9065 16315
rect 400 12430 405 12520
rect 595 12430 600 12520
rect 400 500 600 12430
rect 4925 8655 5025 8660
rect 4925 8565 4930 8655
rect 5020 8565 5025 8655
rect 4925 8560 5025 8565
rect 5415 8655 5515 8660
rect 5415 8565 5420 8655
rect 5510 8565 5515 8655
rect 5415 8560 5515 8565
rect 8475 8655 8575 8660
rect 8475 8565 8480 8655
rect 8570 8565 8575 8655
rect 8475 8560 8575 8565
rect 8965 8655 9065 8660
rect 8965 8565 8970 8655
rect 9060 8565 9065 8655
rect 8965 8560 9065 8565
rect 4950 7285 4980 8560
rect 5435 7530 5465 8560
rect 8510 7685 8540 8560
rect 9005 7860 9035 8560
rect 11385 7860 11415 17650
rect 9005 7830 11415 7860
rect 11605 7685 11635 17930
rect 8510 7655 11635 7685
rect 11865 7530 11895 18180
rect 5435 7500 11895 7530
rect 12195 7285 12225 18425
rect 4910 7255 12225 7285
rect 13250 945 13340 950
rect 13250 855 13255 945
rect 13335 855 13340 945
rect 13250 100 13340 855
rect 15180 620 15270 625
rect 15180 530 15185 620
rect 15265 530 15270 620
rect 15180 100 15270 530
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 100
rect 15181 0 15271 100
use vco  vco_0
timestamp 1725574488
transform 1 0 -970 0 1 10765
box 3265 -3825 12105 6130
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
