magic
tech sky130A
magscale 1 2
timestamp 1725528013
<< pwell >>
rect -367 -686 367 686
<< psubdiff >>
rect -331 616 331 650
rect -331 554 -297 616
rect 297 554 331 616
rect -331 -616 -297 -554
rect 297 -616 331 -554
rect -331 -650 331 -616
<< psubdiffcont >>
rect -331 -554 -297 554
rect 297 -554 331 554
<< xpolycontact >>
rect -201 88 -131 520
rect -201 -520 -131 -88
rect -35 88 35 520
rect -35 -520 35 -88
rect 131 88 201 520
rect 131 -520 201 -88
<< xpolyres >>
rect -201 -88 -131 88
rect -35 -88 35 88
rect 131 -88 201 88
<< locali >>
rect -331 616 331 650
rect -331 554 -297 616
rect 297 554 331 616
rect -331 -616 -297 -554
rect 297 -616 331 -554
rect -331 -650 331 -616
<< viali >>
rect -185 105 -147 502
rect -19 105 19 502
rect 147 105 185 502
rect -185 -502 -147 -105
rect -19 -502 19 -105
rect 147 -502 185 -105
<< metal1 >>
rect -191 502 -141 514
rect -191 105 -185 502
rect -147 105 -141 502
rect -191 93 -141 105
rect -25 502 25 514
rect -25 105 -19 502
rect 19 105 25 502
rect -25 93 25 105
rect 141 502 191 514
rect 141 105 147 502
rect 185 105 191 502
rect 141 93 191 105
rect -191 -105 -141 -93
rect -191 -502 -185 -105
rect -147 -502 -141 -105
rect -191 -514 -141 -502
rect -25 -105 25 -93
rect -25 -502 -19 -105
rect 19 -502 25 -105
rect -25 -514 25 -502
rect 141 -105 191 -93
rect 141 -502 147 -105
rect 185 -502 191 -105
rect 141 -514 191 -502
<< properties >>
string FIXED_BBOX -314 -633 314 633
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.04 m 1 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 7.018k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
