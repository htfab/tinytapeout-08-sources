magic
tech sky130A
magscale 1 2
timestamp 1725572295
<< locali >>
rect 1430 3400 4720 3450
rect 1430 3290 1690 3400
rect 4660 3290 4720 3400
rect 1430 3060 4720 3290
rect 1430 2440 2060 3060
rect 3480 2440 4720 3060
rect 1430 1530 1850 2440
rect 3650 1530 4720 2440
rect 1430 1140 4720 1530
rect 1430 400 2080 1140
rect 3650 1130 4720 1140
rect 4480 400 4720 1130
rect 1430 230 1990 240
rect 1430 -420 4720 230
rect 1430 -2950 1990 -420
rect 4500 -2950 4720 -420
rect 1430 -3380 4720 -2950
rect 1430 -3640 4020 -3380
rect 1430 -3680 2710 -3640
rect 3820 -3680 4020 -3640
rect 1430 -4350 2680 -3680
rect 3850 -4350 4020 -3680
rect 1430 -4490 4020 -4350
rect 1430 -5200 4720 -4490
rect 1430 -5330 1780 -5200
rect 4370 -5330 4720 -5200
rect 1430 -5360 4720 -5330
<< viali >>
rect 1690 3290 4660 3400
rect 1780 -5330 4370 -5200
<< metal1 >>
rect 1430 3400 4720 3450
rect 1430 3290 1690 3400
rect 4660 3290 4720 3400
rect 1430 3250 4720 3290
rect 2010 2900 2020 3100
rect 2230 2900 2240 3100
rect 2010 2290 2020 2490
rect 2220 2290 2230 2490
rect 3300 2290 4330 2490
rect 1430 1640 1630 1710
rect 2010 1700 2020 1900
rect 2220 1700 2230 1900
rect 1430 1570 4720 1640
rect 1430 1510 1630 1570
rect 1430 210 1690 410
rect 1890 350 1900 410
rect 2110 350 2170 980
rect 2370 490 2470 1570
rect 2600 580 2610 980
rect 2680 580 2690 980
rect 2840 500 2940 1570
rect 4370 1400 4570 1460
rect 3470 1320 4570 1400
rect 3120 350 3180 980
rect 3360 350 3420 980
rect 3640 500 3750 1320
rect 3850 580 3860 980
rect 3930 580 3940 980
rect 4090 500 4200 1320
rect 4370 1260 4570 1320
rect 4370 400 4430 980
rect 4370 350 4570 400
rect 1890 270 4570 350
rect 1890 210 1900 270
rect 2070 -2720 2080 -620
rect 2150 -2720 2160 -620
rect 3080 -2860 3310 270
rect 4370 200 4570 270
rect 4340 -2730 4350 -620
rect 4410 -2730 4420 -620
rect 1430 -3040 1630 -3000
rect 4410 -3040 4610 -3000
rect 1430 -3160 4610 -3040
rect 1430 -3200 1630 -3160
rect 2730 -4560 2790 -3780
rect 3000 -4250 3090 -3160
rect 3220 -4180 3230 -3780
rect 3300 -4180 3310 -3780
rect 3450 -4260 3540 -3160
rect 4410 -3200 4610 -3160
rect 3740 -4560 3800 -3780
rect 4520 -4560 4720 -4490
rect 2730 -4620 4720 -4560
rect 4520 -4690 4720 -4620
rect 1430 -5200 4720 -5160
rect 1430 -5330 1780 -5200
rect 4370 -5330 4720 -5200
rect 1430 -5360 4720 -5330
<< via1 >>
rect 1690 3290 4660 3400
rect 2020 2900 2230 3100
rect 2020 2290 2220 2490
rect 2020 1700 2220 1900
rect 1690 210 1890 410
rect 2610 580 2680 980
rect 3860 580 3930 980
rect 2080 -2720 2150 -620
rect 4350 -2730 4410 -620
rect 3230 -4180 3300 -3780
rect 1780 -5330 4370 -5200
<< metal2 >>
rect 1630 3410 3950 3450
rect 1630 3400 4660 3410
rect 1630 3290 1690 3400
rect 1630 3280 4660 3290
rect 1630 3250 3950 3280
rect 2020 3100 2230 3250
rect 2020 2890 2230 2900
rect 2020 2490 2220 2500
rect 2020 2280 2220 2290
rect 2020 1900 2220 1910
rect 2020 1690 2220 1700
rect 1690 410 1890 420
rect 1690 200 1890 210
rect 2090 -610 2150 1690
rect 2620 990 2670 3250
rect 3870 990 3920 3250
rect 2610 980 2680 990
rect 2610 570 2680 580
rect 3860 980 3930 990
rect 3860 570 3930 580
rect 2080 -620 2150 -610
rect 2080 -2730 2150 -2720
rect 2090 -5160 2150 -2730
rect 4350 -620 4410 -580
rect 4350 -3300 4410 -2730
rect 3940 -3360 4410 -3300
rect 3230 -3780 3300 -3770
rect 3230 -4190 3300 -4180
rect 3940 -5160 4000 -3360
rect 1750 -5200 4430 -5160
rect 1750 -5330 1780 -5200
rect 4370 -5330 4430 -5200
rect 1750 -5360 4430 -5330
<< via2 >>
rect 2020 2290 2220 2490
rect 1690 210 1890 410
rect 3230 -4180 3300 -3780
<< metal3 >>
rect 2010 2490 2230 2495
rect 1710 2290 2020 2490
rect 2220 2290 2230 2490
rect 1710 415 1850 2290
rect 2010 2285 2230 2290
rect 1680 410 1900 415
rect 1680 210 1690 410
rect 1890 210 1900 410
rect 1680 205 1900 210
rect 1710 -3930 1850 205
rect 3220 -3780 3310 -3775
rect 3220 -3930 3230 -3780
rect 1710 -4030 3230 -3930
rect 3220 -4180 3230 -4030
rect 3300 -4180 3310 -3780
rect 3220 -4185 3310 -4180
use vco_buffer  vco_buffer_0
timestamp 1725445236
transform 1 0 2020 0 1 1710
box 0 -10 1480 1390
use sky130_fd_pr__nfet_01v8_XVWV9B  XM1
timestamp 1725569918
transform 1 0 3265 0 1 -3980
box -625 -410 625 410
use sky130_fd_pr__pfet_01v8_GJP7VV  XM3
timestamp 1725457726
transform 1 0 2645 0 1 779
box -625 -419 625 419
use sky130_fd_pr__pfet_01v8_GJP7VV  XM7
timestamp 1725457726
transform 1 0 3895 0 1 779
box -625 -419 625 419
use sky130_fd_pr__nfet_01v8_APRB2X  XM8
timestamp 1725457726
transform 1 0 3246 0 1 -1680
box -1296 -1310 1296 1310
<< labels >>
flabel metal1 1430 210 1630 410 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 1430 3250 1630 3450 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 4130 2290 4330 2490 0 FreeSans 256 0 0 0 Vbuf
port 7 nsew
flabel metal1 4370 1260 4570 1460 0 FreeSans 256 0 0 0 Vd
port 4 nsew
flabel metal1 1430 1510 1630 1710 0 FreeSans 256 0 0 0 Vb
port 3 nsew
flabel metal1 1430 -3200 1630 -3000 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 4520 -4690 4720 -4490 0 FreeSans 256 0 0 0 Vs
port 6 nsew
flabel metal1 1430 -5360 1630 -5160 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
