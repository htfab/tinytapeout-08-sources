magic
tech sky130A
magscale 1 2
timestamp 1725172927
<< dnwell >>
rect 10046 10908 12680 12050
<< nwell >>
rect 9966 11844 12760 12130
rect 9966 11114 10252 11844
rect 12474 11114 12760 11844
rect 9966 10828 12760 11114
<< nsubdiff >>
rect 10003 12073 12723 12093
rect 10003 12039 10088 12073
rect 10122 12039 10156 12073
rect 10190 12039 10224 12073
rect 10258 12039 10292 12073
rect 10326 12039 10360 12073
rect 10394 12039 10428 12073
rect 10462 12039 10496 12073
rect 10530 12039 10564 12073
rect 10598 12039 10632 12073
rect 10666 12039 10700 12073
rect 10734 12039 10768 12073
rect 10802 12039 10836 12073
rect 10870 12039 10904 12073
rect 10938 12039 10972 12073
rect 11006 12039 11040 12073
rect 11074 12039 11108 12073
rect 11142 12039 11176 12073
rect 11210 12039 11244 12073
rect 11278 12039 11312 12073
rect 11346 12039 11380 12073
rect 11414 12039 11448 12073
rect 11482 12039 11516 12073
rect 11550 12039 11584 12073
rect 11618 12039 11652 12073
rect 11686 12039 11720 12073
rect 11754 12039 11788 12073
rect 11822 12039 11856 12073
rect 11890 12039 11924 12073
rect 11958 12039 11992 12073
rect 12026 12039 12060 12073
rect 12094 12039 12128 12073
rect 12162 12039 12196 12073
rect 12230 12039 12264 12073
rect 12298 12039 12332 12073
rect 12366 12039 12400 12073
rect 12434 12039 12468 12073
rect 12502 12039 12536 12073
rect 12570 12039 12604 12073
rect 12638 12039 12723 12073
rect 10003 12019 12723 12039
rect 10003 12006 10077 12019
rect 10003 11972 10023 12006
rect 10057 11972 10077 12006
rect 10003 11938 10077 11972
rect 10003 11904 10023 11938
rect 10057 11904 10077 11938
rect 10003 11870 10077 11904
rect 10003 11836 10023 11870
rect 10057 11836 10077 11870
rect 10003 11802 10077 11836
rect 10003 11768 10023 11802
rect 10057 11768 10077 11802
rect 10003 11734 10077 11768
rect 10003 11700 10023 11734
rect 10057 11700 10077 11734
rect 10003 11666 10077 11700
rect 10003 11632 10023 11666
rect 10057 11632 10077 11666
rect 10003 11598 10077 11632
rect 10003 11564 10023 11598
rect 10057 11564 10077 11598
rect 10003 11530 10077 11564
rect 10003 11496 10023 11530
rect 10057 11496 10077 11530
rect 10003 11462 10077 11496
rect 10003 11428 10023 11462
rect 10057 11428 10077 11462
rect 10003 11394 10077 11428
rect 10003 11360 10023 11394
rect 10057 11360 10077 11394
rect 10003 11326 10077 11360
rect 10003 11292 10023 11326
rect 10057 11292 10077 11326
rect 10003 11258 10077 11292
rect 10003 11224 10023 11258
rect 10057 11224 10077 11258
rect 10003 11190 10077 11224
rect 10003 11156 10023 11190
rect 10057 11156 10077 11190
rect 10003 11122 10077 11156
rect 10003 11088 10023 11122
rect 10057 11088 10077 11122
rect 10003 11054 10077 11088
rect 10003 11020 10023 11054
rect 10057 11020 10077 11054
rect 10003 10986 10077 11020
rect 10003 10952 10023 10986
rect 10057 10952 10077 10986
rect 10003 10939 10077 10952
rect 12649 12006 12723 12019
rect 12649 11972 12669 12006
rect 12703 11972 12723 12006
rect 12649 11938 12723 11972
rect 12649 11904 12669 11938
rect 12703 11904 12723 11938
rect 12649 11870 12723 11904
rect 12649 11836 12669 11870
rect 12703 11836 12723 11870
rect 12649 11802 12723 11836
rect 12649 11768 12669 11802
rect 12703 11768 12723 11802
rect 12649 11734 12723 11768
rect 12649 11700 12669 11734
rect 12703 11700 12723 11734
rect 12649 11666 12723 11700
rect 12649 11632 12669 11666
rect 12703 11632 12723 11666
rect 12649 11598 12723 11632
rect 12649 11564 12669 11598
rect 12703 11564 12723 11598
rect 12649 11530 12723 11564
rect 12649 11496 12669 11530
rect 12703 11496 12723 11530
rect 12649 11462 12723 11496
rect 12649 11428 12669 11462
rect 12703 11428 12723 11462
rect 12649 11394 12723 11428
rect 12649 11360 12669 11394
rect 12703 11360 12723 11394
rect 12649 11326 12723 11360
rect 12649 11292 12669 11326
rect 12703 11292 12723 11326
rect 12649 11258 12723 11292
rect 12649 11224 12669 11258
rect 12703 11224 12723 11258
rect 12649 11190 12723 11224
rect 12649 11156 12669 11190
rect 12703 11156 12723 11190
rect 12649 11122 12723 11156
rect 12649 11088 12669 11122
rect 12703 11088 12723 11122
rect 12649 11054 12723 11088
rect 12649 11020 12669 11054
rect 12703 11020 12723 11054
rect 12649 10986 12723 11020
rect 12649 10952 12669 10986
rect 12703 10952 12723 10986
rect 12649 10939 12723 10952
rect 10003 10919 12723 10939
rect 10003 10885 10088 10919
rect 10122 10885 10156 10919
rect 10190 10885 10224 10919
rect 10258 10885 10292 10919
rect 10326 10885 10360 10919
rect 10394 10885 10428 10919
rect 10462 10885 10496 10919
rect 10530 10885 10564 10919
rect 10598 10885 10632 10919
rect 10666 10885 10700 10919
rect 10734 10885 10768 10919
rect 10802 10885 10836 10919
rect 10870 10885 10904 10919
rect 10938 10885 10972 10919
rect 11006 10885 11040 10919
rect 11074 10885 11108 10919
rect 11142 10885 11176 10919
rect 11210 10885 11244 10919
rect 11278 10885 11312 10919
rect 11346 10885 11380 10919
rect 11414 10885 11448 10919
rect 11482 10885 11516 10919
rect 11550 10885 11584 10919
rect 11618 10885 11652 10919
rect 11686 10885 11720 10919
rect 11754 10885 11788 10919
rect 11822 10885 11856 10919
rect 11890 10885 11924 10919
rect 11958 10885 11992 10919
rect 12026 10885 12060 10919
rect 12094 10885 12128 10919
rect 12162 10885 12196 10919
rect 12230 10885 12264 10919
rect 12298 10885 12332 10919
rect 12366 10885 12400 10919
rect 12434 10885 12468 10919
rect 12502 10885 12536 10919
rect 12570 10885 12604 10919
rect 12638 10885 12723 10919
rect 10003 10865 12723 10885
<< nsubdiffcont >>
rect 10088 12039 10122 12073
rect 10156 12039 10190 12073
rect 10224 12039 10258 12073
rect 10292 12039 10326 12073
rect 10360 12039 10394 12073
rect 10428 12039 10462 12073
rect 10496 12039 10530 12073
rect 10564 12039 10598 12073
rect 10632 12039 10666 12073
rect 10700 12039 10734 12073
rect 10768 12039 10802 12073
rect 10836 12039 10870 12073
rect 10904 12039 10938 12073
rect 10972 12039 11006 12073
rect 11040 12039 11074 12073
rect 11108 12039 11142 12073
rect 11176 12039 11210 12073
rect 11244 12039 11278 12073
rect 11312 12039 11346 12073
rect 11380 12039 11414 12073
rect 11448 12039 11482 12073
rect 11516 12039 11550 12073
rect 11584 12039 11618 12073
rect 11652 12039 11686 12073
rect 11720 12039 11754 12073
rect 11788 12039 11822 12073
rect 11856 12039 11890 12073
rect 11924 12039 11958 12073
rect 11992 12039 12026 12073
rect 12060 12039 12094 12073
rect 12128 12039 12162 12073
rect 12196 12039 12230 12073
rect 12264 12039 12298 12073
rect 12332 12039 12366 12073
rect 12400 12039 12434 12073
rect 12468 12039 12502 12073
rect 12536 12039 12570 12073
rect 12604 12039 12638 12073
rect 10023 11972 10057 12006
rect 10023 11904 10057 11938
rect 10023 11836 10057 11870
rect 10023 11768 10057 11802
rect 10023 11700 10057 11734
rect 10023 11632 10057 11666
rect 10023 11564 10057 11598
rect 10023 11496 10057 11530
rect 10023 11428 10057 11462
rect 10023 11360 10057 11394
rect 10023 11292 10057 11326
rect 10023 11224 10057 11258
rect 10023 11156 10057 11190
rect 10023 11088 10057 11122
rect 10023 11020 10057 11054
rect 10023 10952 10057 10986
rect 12669 11972 12703 12006
rect 12669 11904 12703 11938
rect 12669 11836 12703 11870
rect 12669 11768 12703 11802
rect 12669 11700 12703 11734
rect 12669 11632 12703 11666
rect 12669 11564 12703 11598
rect 12669 11496 12703 11530
rect 12669 11428 12703 11462
rect 12669 11360 12703 11394
rect 12669 11292 12703 11326
rect 12669 11224 12703 11258
rect 12669 11156 12703 11190
rect 12669 11088 12703 11122
rect 12669 11020 12703 11054
rect 12669 10952 12703 10986
rect 10088 10885 10122 10919
rect 10156 10885 10190 10919
rect 10224 10885 10258 10919
rect 10292 10885 10326 10919
rect 10360 10885 10394 10919
rect 10428 10885 10462 10919
rect 10496 10885 10530 10919
rect 10564 10885 10598 10919
rect 10632 10885 10666 10919
rect 10700 10885 10734 10919
rect 10768 10885 10802 10919
rect 10836 10885 10870 10919
rect 10904 10885 10938 10919
rect 10972 10885 11006 10919
rect 11040 10885 11074 10919
rect 11108 10885 11142 10919
rect 11176 10885 11210 10919
rect 11244 10885 11278 10919
rect 11312 10885 11346 10919
rect 11380 10885 11414 10919
rect 11448 10885 11482 10919
rect 11516 10885 11550 10919
rect 11584 10885 11618 10919
rect 11652 10885 11686 10919
rect 11720 10885 11754 10919
rect 11788 10885 11822 10919
rect 11856 10885 11890 10919
rect 11924 10885 11958 10919
rect 11992 10885 12026 10919
rect 12060 10885 12094 10919
rect 12128 10885 12162 10919
rect 12196 10885 12230 10919
rect 12264 10885 12298 10919
rect 12332 10885 12366 10919
rect 12400 10885 12434 10919
rect 12468 10885 12502 10919
rect 12536 10885 12570 10919
rect 12604 10885 12638 10919
<< locali >>
rect 10023 12039 10088 12073
rect 10122 12039 10156 12073
rect 10190 12039 10224 12073
rect 10258 12039 10292 12073
rect 10326 12039 10360 12073
rect 10394 12039 10428 12073
rect 10462 12039 10496 12073
rect 10530 12039 10564 12073
rect 10598 12039 10632 12073
rect 10666 12039 10700 12073
rect 10734 12039 10768 12073
rect 10802 12039 10836 12073
rect 10870 12039 10904 12073
rect 10938 12039 10972 12073
rect 11006 12039 11040 12073
rect 11074 12039 11108 12073
rect 11142 12039 11176 12073
rect 11210 12039 11244 12073
rect 11278 12039 11312 12073
rect 11346 12039 11380 12073
rect 11414 12039 11448 12073
rect 11482 12039 11516 12073
rect 11550 12039 11584 12073
rect 11618 12039 11652 12073
rect 11686 12039 11720 12073
rect 11754 12039 11788 12073
rect 11822 12039 11856 12073
rect 11890 12039 11924 12073
rect 11958 12039 11992 12073
rect 12026 12039 12060 12073
rect 12094 12039 12128 12073
rect 12162 12039 12196 12073
rect 12230 12039 12264 12073
rect 12298 12039 12332 12073
rect 12366 12039 12400 12073
rect 12434 12039 12468 12073
rect 12502 12039 12536 12073
rect 12570 12039 12604 12073
rect 12638 12039 12703 12073
rect 10023 12006 10057 12039
rect 10023 11938 10057 11972
rect 10023 11870 10057 11904
rect 10023 11802 10057 11836
rect 10023 11734 10057 11768
rect 10023 11666 10057 11700
rect 10023 11598 10057 11632
rect 12669 12006 12703 12039
rect 12669 11938 12703 11972
rect 12669 11870 12703 11904
rect 12669 11802 12703 11836
rect 12669 11734 12703 11768
rect 12669 11666 12703 11700
rect 12669 11598 12703 11632
rect 10023 11530 10057 11564
rect 12302 11500 12350 11568
rect 12669 11530 12703 11564
rect 10023 11462 10057 11496
rect 10023 11394 10057 11428
rect 10023 11326 10057 11360
rect 10023 11258 10057 11292
rect 10023 11190 10057 11224
rect 12669 11462 12703 11496
rect 12669 11394 12703 11428
rect 12669 11326 12703 11360
rect 12669 11258 12703 11292
rect 10023 11122 10057 11156
rect 10023 11054 10057 11088
rect 10023 10986 10057 11020
rect 11840 11176 12110 11196
rect 11840 10998 11850 11176
rect 12100 10998 12110 11176
rect 11840 10978 12110 10998
rect 12669 11190 12703 11224
rect 12669 11122 12703 11156
rect 12669 11054 12703 11088
rect 12669 10986 12703 11020
rect 10023 10919 10057 10952
rect 12669 10919 12703 10952
rect 10023 10885 10088 10919
rect 10122 10885 10156 10919
rect 10190 10885 10224 10919
rect 10258 10885 10292 10919
rect 10326 10885 10360 10919
rect 10394 10885 10428 10919
rect 10462 10885 10496 10919
rect 10530 10885 10564 10919
rect 10598 10885 10632 10919
rect 10666 10885 10700 10919
rect 10734 10885 10768 10919
rect 10802 10885 10836 10919
rect 10870 10885 10904 10919
rect 10938 10885 10972 10919
rect 11006 10885 11040 10919
rect 11074 10885 11108 10919
rect 11142 10885 11176 10919
rect 11210 10885 11244 10919
rect 11278 10885 11312 10919
rect 11346 10885 11380 10919
rect 11414 10885 11448 10919
rect 11482 10885 11516 10919
rect 11550 10885 11584 10919
rect 11618 10885 11652 10919
rect 11686 10885 11720 10919
rect 11754 10885 11788 10919
rect 11822 10885 11856 10919
rect 11890 10885 11924 10919
rect 11958 10885 11992 10919
rect 12026 10885 12060 10919
rect 12094 10885 12128 10919
rect 12162 10885 12196 10919
rect 12230 10885 12264 10919
rect 12298 10885 12332 10919
rect 12366 10885 12400 10919
rect 12434 10885 12468 10919
rect 12502 10885 12536 10919
rect 12570 10885 12604 10919
rect 12638 10885 12703 10919
rect 6568 10108 6718 10170
rect 4138 9548 4732 9696
rect 10356 9686 10406 9706
rect 10356 9652 10364 9686
rect 10398 9652 10406 9686
rect 10356 9614 10406 9652
rect 10356 9580 10364 9614
rect 10398 9580 10406 9614
rect 10356 9560 10406 9580
rect 4142 5642 4298 9548
rect 6590 9056 6736 9130
rect 8098 8929 8148 8958
rect 8098 8895 8106 8929
rect 8140 8895 8148 8929
rect 8098 8866 8148 8895
rect 11982 8758 14642 8900
rect 8114 8362 8514 8384
rect 8672 8362 8698 8384
rect 7878 8285 7948 8286
rect 7878 8251 7896 8285
rect 7930 8251 7948 8285
rect 8114 8260 8698 8362
rect 7878 8213 7948 8251
rect 7878 8179 7896 8213
rect 7930 8179 7948 8213
rect 7878 8178 7948 8179
rect 6614 7942 6760 8016
rect 14326 7808 14420 7884
rect 8008 7582 8068 7630
rect 6314 7124 6372 7172
rect 11280 7146 11336 7150
rect 8062 6968 8222 7142
rect 11280 7112 11291 7146
rect 11325 7112 11336 7146
rect 11280 7108 11336 7112
rect 10918 7086 10954 7088
rect 10918 7052 10919 7086
rect 10953 7052 10954 7086
rect 10918 7050 10954 7052
rect 11084 7017 11146 7024
rect 11084 6983 11098 7017
rect 11132 6983 11146 7017
rect 11084 6976 11146 6983
rect 10010 6941 10066 6946
rect 10010 6907 10021 6941
rect 10055 6907 10066 6941
rect 10010 6904 10066 6907
rect 8500 6532 8634 6850
rect 14540 6766 14636 8758
rect 11506 6714 14642 6766
rect 11344 6678 14642 6714
rect 10344 6516 10484 6518
rect 10344 6482 10361 6516
rect 10395 6482 10433 6516
rect 10467 6482 10484 6516
rect 10344 6480 10484 6482
rect 7792 6144 7944 6218
rect 4596 5642 4710 6002
rect 4142 5534 4710 5642
rect 5442 5821 5552 5838
rect 5442 5643 5444 5821
rect 5550 5643 5552 5821
rect 8706 5774 9052 5884
rect 8426 5702 8484 5750
rect 9028 5709 9206 5724
rect 9062 5675 9100 5709
rect 9134 5675 9172 5709
rect 9028 5660 9206 5675
rect 5442 5626 5552 5643
rect 4148 5526 4710 5534
rect 4430 4777 4486 4780
rect 4288 4774 4330 4776
rect 4288 4740 4292 4774
rect 4326 4740 4330 4774
rect 4430 4743 4441 4777
rect 4475 4743 4486 4777
rect 4430 4740 4486 4743
rect 4288 4738 4330 4740
rect 4596 4676 4710 5526
rect 6410 5396 6468 5444
rect 4596 4570 5878 4676
rect 4596 4538 4710 4570
rect 4458 4502 4710 4538
<< viali >>
rect 11850 10998 12100 11176
rect 10364 9652 10398 9686
rect 10364 9580 10398 9614
rect 8106 8895 8140 8929
rect 7896 8251 7930 8285
rect 7896 8179 7930 8213
rect 11291 7112 11325 7146
rect 10919 7052 10953 7086
rect 10122 6978 10156 7012
rect 11098 6983 11132 7017
rect 10021 6907 10055 6941
rect 10361 6482 10395 6516
rect 10433 6482 10467 6516
rect 5444 5643 5550 5821
rect 9028 5675 9062 5709
rect 9100 5675 9134 5709
rect 9172 5675 9206 5709
rect 4292 4740 4326 4774
rect 4441 4743 4475 4777
<< metal1 >>
rect 8272 11936 8530 11958
rect 8257 11934 12358 11936
rect 8257 11814 12360 11934
rect 6772 10919 7008 10936
rect 6772 10739 6800 10919
rect 6980 10739 7008 10919
rect 6772 10722 7008 10739
rect 7602 10682 8112 10698
rect 8272 10682 8530 11814
rect 10368 11662 10432 11814
rect 10368 11406 10434 11662
rect 10684 11656 10711 11708
rect 10763 11656 10775 11708
rect 10827 11656 10839 11708
rect 10891 11656 10903 11708
rect 10955 11656 10967 11708
rect 11019 11656 11031 11708
rect 11083 11656 11095 11708
rect 11147 11656 11159 11708
rect 11211 11656 11223 11708
rect 11275 11656 11287 11708
rect 11339 11656 11351 11708
rect 11403 11656 11415 11708
rect 11467 11656 11479 11708
rect 11531 11656 11558 11708
rect 11724 11607 12200 11608
rect 11724 11555 11744 11607
rect 11796 11555 11808 11607
rect 11860 11555 11872 11607
rect 11924 11555 11936 11607
rect 11988 11555 12000 11607
rect 12052 11555 12064 11607
rect 12116 11555 12128 11607
rect 12180 11555 12200 11607
rect 12306 11566 12360 11814
rect 11724 11554 12200 11555
rect 10688 11462 10715 11514
rect 10767 11462 10779 11514
rect 10831 11462 10843 11514
rect 10895 11462 10907 11514
rect 10959 11462 10971 11514
rect 11023 11462 11035 11514
rect 11087 11462 11099 11514
rect 11151 11462 11163 11514
rect 11215 11462 11227 11514
rect 11279 11462 11291 11514
rect 11343 11462 11355 11514
rect 11407 11462 11419 11514
rect 11471 11462 11483 11514
rect 11535 11462 11562 11514
rect 10370 11404 10434 11406
rect 11716 11419 12192 11420
rect 11716 11367 11736 11419
rect 11788 11367 11800 11419
rect 11852 11367 11864 11419
rect 11916 11367 11928 11419
rect 11980 11367 11992 11419
rect 12044 11367 12056 11419
rect 12108 11367 12120 11419
rect 12172 11367 12192 11419
rect 11716 11366 12192 11367
rect 10698 11262 10725 11314
rect 10777 11262 10789 11314
rect 10841 11262 10853 11314
rect 10905 11262 10917 11314
rect 10969 11262 10981 11314
rect 11033 11262 11045 11314
rect 11097 11262 11109 11314
rect 11161 11262 11173 11314
rect 11225 11262 11237 11314
rect 11289 11262 11301 11314
rect 11353 11262 11365 11314
rect 11417 11262 11429 11314
rect 11481 11262 11493 11314
rect 11545 11262 11572 11314
rect 12296 11308 12360 11566
rect 12296 11306 12352 11308
rect 11828 11177 12122 11202
rect 11828 11176 11853 11177
rect 12097 11176 12122 11177
rect 7602 10596 8530 10682
rect 8924 11058 8980 11078
rect 11828 11058 11850 11176
rect 8924 10998 11850 11058
rect 12100 10998 12122 11176
rect 8924 10997 11853 10998
rect 12097 10997 12122 10998
rect 8924 10972 12122 10997
rect 8924 10936 12098 10972
rect 7602 10590 8448 10596
rect 7602 10570 8112 10590
rect 5544 10482 6562 10496
rect 5484 10408 6562 10482
rect 5484 10378 5550 10408
rect 5484 10365 5566 10378
rect 4830 10325 5108 10346
rect 4830 9953 4847 10325
rect 5091 9953 5108 10325
rect 4830 9932 5108 9953
rect 5484 10313 5499 10365
rect 5551 10313 5566 10365
rect 5484 10301 5566 10313
rect 5484 10249 5499 10301
rect 5551 10249 5566 10301
rect 5484 10237 5566 10249
rect 5484 10185 5499 10237
rect 5551 10185 5566 10237
rect 5484 10173 5566 10185
rect 5484 10121 5499 10173
rect 5551 10121 5566 10173
rect 5484 10109 5566 10121
rect 5484 10057 5499 10109
rect 5551 10057 5566 10109
rect 5484 10045 5566 10057
rect 5484 9993 5499 10045
rect 5551 9993 5566 10045
rect 5484 9980 5566 9993
rect 6550 10367 6624 10378
rect 6550 10315 6561 10367
rect 6613 10315 6624 10367
rect 6550 10303 6624 10315
rect 6550 10251 6561 10303
rect 6613 10251 6624 10303
rect 6550 10239 6624 10251
rect 6550 10187 6561 10239
rect 6613 10187 6624 10239
rect 6550 10175 6624 10187
rect 6550 10123 6561 10175
rect 6613 10123 6624 10175
rect 6550 10111 6624 10123
rect 6662 10249 6742 10262
rect 6662 10197 6676 10249
rect 6728 10197 6742 10249
rect 6662 10185 6742 10197
rect 6662 10133 6676 10185
rect 6728 10133 6742 10185
rect 6662 10120 6742 10133
rect 6550 10059 6561 10111
rect 6613 10059 6624 10111
rect 6550 10047 6624 10059
rect 6550 9995 6561 10047
rect 6613 9995 6624 10047
rect 6550 9984 6624 9995
rect 7576 10004 7648 10024
rect 5484 9950 5550 9980
rect 7576 9952 7586 10004
rect 7638 9952 7648 10004
rect 5484 9862 6602 9950
rect 7576 9940 7648 9952
rect 7576 9888 7586 9940
rect 7638 9888 7648 9940
rect 7576 9868 7648 9888
rect 7778 10002 7850 10022
rect 7778 9950 7788 10002
rect 7840 9950 7850 10002
rect 7778 9938 7850 9950
rect 7778 9886 7788 9938
rect 7840 9886 7850 9938
rect 7778 9866 7850 9886
rect 7966 10008 8038 10028
rect 7966 9956 7976 10008
rect 8028 9956 8038 10008
rect 7966 9944 8038 9956
rect 7966 9892 7976 9944
rect 8028 9892 8038 9944
rect 7966 9872 8038 9892
rect 4826 9687 5104 9708
rect 4826 9682 4843 9687
rect 4794 9315 4843 9682
rect 5087 9315 5104 9687
rect 5886 9692 6136 9862
rect 6832 9692 6930 9698
rect 5886 9592 6938 9692
rect 5510 9392 5592 9398
rect 5508 9316 6576 9392
rect 4794 9294 5104 9315
rect 4346 8764 4574 8780
rect 4794 8764 5088 9294
rect 5510 9244 5592 9316
rect 5506 9213 5592 9244
rect 5506 9161 5517 9213
rect 5569 9161 5592 9213
rect 6832 9180 6930 9592
rect 5506 9149 5592 9161
rect 5506 9097 5517 9149
rect 5569 9097 5592 9149
rect 5506 9085 5592 9097
rect 5506 9033 5517 9085
rect 5569 9033 5592 9085
rect 5506 9002 5592 9033
rect 5510 8856 5592 9002
rect 6558 9179 6978 9180
rect 6558 9127 6581 9179
rect 6633 9156 6978 9179
rect 6633 9127 6703 9156
rect 6558 9115 6703 9127
rect 6558 9063 6581 9115
rect 6633 9104 6703 9115
rect 6755 9104 6978 9156
rect 6633 9092 6978 9104
rect 6633 9063 6703 9092
rect 6558 9051 6703 9063
rect 6558 8999 6581 9051
rect 6633 9040 6703 9051
rect 6755 9040 6978 9092
rect 6633 8999 6978 9040
rect 6558 8998 6978 8999
rect 6574 8996 6978 8998
rect 6832 8992 6930 8996
rect 7676 8970 7748 8990
rect 7676 8918 7686 8970
rect 7738 8918 7748 8970
rect 7676 8906 7748 8918
rect 5950 8856 6146 8874
rect 5510 8792 6578 8856
rect 7676 8854 7686 8906
rect 7738 8854 7748 8906
rect 7676 8834 7748 8854
rect 7874 8964 7946 8984
rect 8092 8966 8154 8970
rect 7874 8912 7884 8964
rect 7936 8912 7946 8964
rect 7874 8900 7946 8912
rect 7874 8848 7884 8900
rect 7936 8848 7946 8900
rect 8088 8945 8164 8966
rect 8088 8893 8100 8945
rect 8152 8893 8164 8945
rect 8088 8872 8164 8893
rect 8092 8854 8154 8872
rect 7874 8828 7946 8848
rect 5510 8766 5592 8792
rect 4346 8552 5088 8764
rect 5950 8730 6146 8792
rect 5954 8604 6144 8730
rect 7494 8706 8004 8708
rect 8256 8706 8336 10590
rect 7494 8620 8646 8706
rect 6862 8604 6972 8606
rect 4346 7726 4574 8552
rect 4794 8550 5088 8552
rect 5946 8518 6972 8604
rect 7494 8580 8004 8620
rect 6062 8516 6972 8518
rect 5542 8274 5606 8276
rect 5542 8206 6600 8274
rect 5542 8174 5606 8206
rect 5528 8161 5610 8174
rect 5528 8109 5543 8161
rect 5595 8109 5610 8161
rect 5528 8097 5610 8109
rect 5528 8045 5543 8097
rect 5595 8045 5610 8097
rect 5528 8033 5610 8045
rect 5528 7981 5543 8033
rect 5595 7981 5610 8033
rect 5528 7969 5610 7981
rect 5528 7917 5543 7969
rect 5595 7917 5610 7969
rect 5528 7905 5610 7917
rect 5528 7853 5543 7905
rect 5595 7853 5610 7905
rect 6588 8100 6698 8178
rect 6588 8098 6694 8100
rect 6588 8046 6606 8098
rect 6658 8052 6694 8098
rect 6862 8052 6972 8516
rect 6658 8046 6972 8052
rect 6588 8034 6730 8046
rect 6588 7982 6606 8034
rect 6658 7994 6730 8034
rect 6782 7994 6972 8046
rect 6658 7982 6972 7994
rect 6588 7970 6730 7982
rect 6588 7918 6606 7970
rect 6658 7930 6730 7970
rect 6782 7930 6972 7982
rect 6658 7922 6972 7930
rect 6658 7918 6694 7922
rect 6588 7900 6694 7918
rect 5528 7841 5610 7853
rect 5528 7789 5543 7841
rect 5595 7789 5610 7841
rect 5528 7776 5610 7789
rect 6584 7782 6690 7900
rect 5542 7736 5606 7776
rect 5160 7732 5654 7736
rect 5160 7728 6592 7732
rect 4346 7719 4900 7726
rect 4346 7539 4371 7719
rect 4551 7539 4900 7719
rect 4346 7528 4900 7539
rect 4354 7526 4900 7528
rect 4636 7158 4900 7526
rect 5154 7678 6592 7728
rect 5154 7662 5654 7678
rect 7564 7676 7818 8580
rect 7872 8286 7954 8298
rect 7994 8288 8056 8338
rect 7868 8285 7958 8286
rect 7868 8258 7896 8285
rect 7930 8258 7958 8285
rect 7868 8206 7887 8258
rect 7939 8206 7958 8258
rect 7994 8210 8068 8288
rect 8728 8210 8778 8296
rect 7994 8208 8802 8210
rect 8924 8208 8980 10936
rect 9352 10506 9538 10510
rect 9232 10488 9638 10506
rect 9232 10308 9249 10488
rect 9621 10308 9638 10488
rect 9232 10290 9638 10308
rect 9352 9814 9538 10290
rect 11616 9841 11884 9866
rect 9352 9812 9864 9814
rect 9352 9740 10284 9812
rect 9352 9738 9864 9740
rect 9352 9276 9538 9738
rect 10350 9686 10412 9718
rect 9728 9646 9822 9672
rect 9728 9594 9749 9646
rect 9801 9594 9822 9646
rect 9728 9568 9822 9594
rect 9936 9640 10010 9666
rect 9936 9588 9947 9640
rect 9999 9588 10010 9640
rect 9936 9562 10010 9588
rect 10122 9638 10196 9664
rect 10350 9660 10364 9686
rect 10122 9586 10133 9638
rect 10185 9586 10196 9638
rect 10122 9560 10196 9586
rect 10346 9652 10364 9660
rect 10398 9660 10412 9686
rect 10398 9652 10434 9660
rect 10346 9636 10434 9652
rect 10346 9580 10364 9636
rect 10416 9584 10434 9636
rect 10398 9580 10434 9584
rect 10346 9560 10434 9580
rect 10350 9548 10412 9560
rect 11616 9469 11628 9841
rect 11872 9469 11884 9841
rect 11616 9444 11884 9469
rect 9838 9410 9912 9436
rect 9838 9358 9849 9410
rect 9901 9358 9912 9410
rect 9838 9332 9912 9358
rect 10028 9408 10102 9434
rect 10028 9356 10039 9408
rect 10091 9356 10102 9408
rect 10028 9330 10102 9356
rect 10220 9412 10294 9438
rect 10220 9360 10231 9412
rect 10283 9360 10294 9412
rect 10220 9334 10294 9360
rect 9352 9274 9986 9276
rect 9352 9202 10276 9274
rect 9352 9190 9986 9202
rect 9490 9186 9986 9190
rect 11596 9201 11898 9218
rect 11596 8829 11625 9201
rect 11869 8829 11898 9201
rect 11596 8812 11898 8829
rect 7868 8179 7896 8206
rect 7930 8179 7958 8206
rect 7868 8178 7958 8179
rect 7996 8199 9022 8208
rect 7872 8166 7954 8178
rect 7996 8160 8358 8199
rect 8008 8154 8358 8160
rect 8338 8147 8358 8154
rect 8410 8147 8422 8199
rect 8474 8162 9022 8199
rect 8474 8154 8802 8162
rect 8924 8158 8980 8162
rect 8474 8147 8494 8154
rect 8338 8146 8494 8147
rect 9206 7957 9288 7972
rect 9206 7905 9221 7957
rect 9273 7905 9288 7957
rect 9206 7893 9288 7905
rect 9206 7841 9221 7893
rect 9273 7841 9288 7893
rect 9206 7829 9288 7841
rect 9206 7777 9221 7829
rect 9273 7777 9288 7829
rect 14276 7961 14348 7964
rect 14276 7909 14286 7961
rect 14338 7909 14348 7961
rect 14276 7897 14348 7909
rect 14276 7845 14286 7897
rect 14338 7845 14348 7897
rect 14276 7833 14348 7845
rect 14276 7781 14286 7833
rect 14338 7781 14348 7833
rect 14276 7778 14348 7781
rect 9206 7762 9288 7777
rect 7558 7670 8570 7676
rect 4616 7127 4912 7158
rect 4616 6755 4642 7127
rect 4886 6755 4912 7127
rect 4616 6724 4912 6755
rect 4636 6722 4900 6724
rect 4616 6457 4912 6488
rect 4078 6402 4544 6404
rect 4616 6402 4642 6457
rect 3574 6398 3848 6400
rect 4078 6398 4642 6402
rect 3574 6116 4642 6398
rect 3574 6110 4110 6116
rect 4458 6110 4642 6116
rect 3574 4788 3848 6110
rect 4616 6085 4642 6110
rect 4886 6402 4912 6457
rect 4886 6110 4924 6402
rect 4886 6085 4912 6110
rect 4616 6054 4912 6085
rect 5154 5842 5334 7662
rect 7548 7570 8570 7670
rect 7548 7530 7802 7570
rect 7548 7408 7818 7530
rect 8462 7492 8564 7570
rect 7564 7268 7818 7408
rect 7916 7417 8030 7438
rect 8462 7424 9092 7492
rect 8468 7420 9092 7424
rect 7916 7365 7947 7417
rect 7999 7365 8030 7417
rect 7916 7353 8030 7365
rect 7916 7301 7947 7353
rect 7999 7301 8030 7353
rect 7916 7280 8030 7301
rect 8398 7351 8474 7378
rect 8398 7299 8410 7351
rect 8462 7299 8474 7351
rect 8398 7272 8474 7299
rect 8590 7349 8666 7376
rect 8590 7297 8602 7349
rect 8654 7297 8666 7349
rect 8590 7270 8666 7297
rect 8792 7347 8868 7374
rect 8792 7295 8804 7347
rect 8856 7295 8868 7347
rect 8792 7268 8868 7295
rect 6500 7194 6968 7228
rect 5732 7112 6968 7194
rect 5582 7070 5660 7080
rect 5582 7018 5595 7070
rect 5647 7018 5660 7070
rect 5582 7006 5660 7018
rect 5582 6954 5595 7006
rect 5647 6954 5660 7006
rect 5582 6942 5660 6954
rect 5582 6890 5595 6942
rect 5647 6890 5660 6942
rect 5582 6878 5660 6890
rect 5582 6826 5595 6878
rect 5647 6826 5660 6878
rect 5582 6814 5660 6826
rect 5582 6762 5595 6814
rect 5647 6762 5660 6814
rect 5582 6750 5660 6762
rect 5582 6698 5595 6750
rect 5647 6698 5660 6750
rect 5582 6686 5660 6698
rect 5582 6634 5595 6686
rect 5647 6634 5660 6686
rect 5582 6624 5660 6634
rect 5774 7066 5852 7076
rect 5774 7014 5787 7066
rect 5839 7014 5852 7066
rect 5774 7002 5852 7014
rect 5774 6950 5787 7002
rect 5839 6950 5852 7002
rect 5774 6938 5852 6950
rect 5774 6886 5787 6938
rect 5839 6886 5852 6938
rect 5774 6874 5852 6886
rect 5774 6822 5787 6874
rect 5839 6822 5852 6874
rect 5774 6810 5852 6822
rect 5774 6758 5787 6810
rect 5839 6758 5852 6810
rect 5774 6746 5852 6758
rect 5774 6694 5787 6746
rect 5839 6694 5852 6746
rect 5774 6682 5852 6694
rect 5774 6630 5787 6682
rect 5839 6630 5852 6682
rect 5774 6620 5852 6630
rect 5968 7072 6046 7082
rect 5968 7020 5981 7072
rect 6033 7020 6046 7072
rect 5968 7008 6046 7020
rect 5968 6956 5981 7008
rect 6033 6956 6046 7008
rect 5968 6944 6046 6956
rect 5968 6892 5981 6944
rect 6033 6892 6046 6944
rect 5968 6880 6046 6892
rect 5968 6828 5981 6880
rect 6033 6828 6046 6880
rect 5968 6816 6046 6828
rect 5968 6764 5981 6816
rect 6033 6764 6046 6816
rect 5968 6752 6046 6764
rect 5968 6700 5981 6752
rect 6033 6700 6046 6752
rect 5968 6688 6046 6700
rect 5968 6636 5981 6688
rect 6033 6636 6046 6688
rect 5968 6626 6046 6636
rect 6160 7070 6238 7080
rect 6160 7018 6173 7070
rect 6225 7018 6238 7070
rect 6160 7006 6238 7018
rect 6160 6954 6173 7006
rect 6225 6954 6238 7006
rect 6160 6942 6238 6954
rect 6160 6890 6173 6942
rect 6225 6890 6238 6942
rect 6160 6878 6238 6890
rect 6160 6826 6173 6878
rect 6225 6826 6238 6878
rect 6160 6814 6238 6826
rect 6160 6762 6173 6814
rect 6225 6762 6238 6814
rect 6160 6750 6238 6762
rect 6160 6698 6173 6750
rect 6225 6698 6238 6750
rect 6160 6686 6238 6698
rect 6160 6634 6173 6686
rect 6225 6634 6238 6686
rect 6160 6624 6238 6634
rect 6354 7070 6432 7080
rect 6354 7018 6367 7070
rect 6419 7018 6432 7070
rect 6354 7006 6432 7018
rect 6354 6954 6367 7006
rect 6419 6954 6432 7006
rect 6354 6942 6432 6954
rect 6354 6890 6367 6942
rect 6419 6890 6432 6942
rect 6354 6878 6432 6890
rect 6354 6826 6367 6878
rect 6419 6826 6432 6878
rect 6354 6814 6432 6826
rect 6354 6762 6367 6814
rect 6419 6762 6432 6814
rect 6354 6750 6432 6762
rect 6354 6698 6367 6750
rect 6419 6698 6432 6750
rect 6354 6686 6432 6698
rect 6354 6634 6367 6686
rect 6419 6634 6432 6686
rect 6354 6624 6432 6634
rect 6546 7066 6624 7076
rect 6546 7014 6559 7066
rect 6611 7014 6624 7066
rect 6546 7002 6624 7014
rect 6546 6950 6559 7002
rect 6611 6950 6624 7002
rect 6546 6938 6624 6950
rect 6546 6886 6559 6938
rect 6611 6886 6624 6938
rect 6546 6874 6624 6886
rect 6546 6822 6559 6874
rect 6611 6822 6624 6874
rect 6546 6810 6624 6822
rect 6546 6758 6559 6810
rect 6611 6758 6624 6810
rect 6546 6746 6624 6758
rect 6546 6694 6559 6746
rect 6611 6694 6624 6746
rect 6546 6682 6624 6694
rect 6546 6630 6559 6682
rect 6611 6630 6624 6682
rect 6546 6620 6624 6630
rect 5872 5966 5950 5976
rect 5678 5962 5756 5966
rect 5678 5910 5691 5962
rect 5743 5910 5756 5962
rect 5678 5898 5756 5910
rect 5160 5834 5362 5842
rect 5436 5834 5558 5850
rect 5678 5846 5691 5898
rect 5743 5846 5756 5898
rect 5678 5834 5756 5846
rect 5872 5914 5885 5966
rect 5937 5914 5950 5966
rect 5872 5902 5950 5914
rect 5872 5850 5885 5902
rect 5937 5850 5950 5902
rect 5872 5838 5950 5850
rect 5160 5832 5558 5834
rect 5160 5821 5473 5832
rect 5525 5821 5558 5832
rect 5160 5650 5444 5821
rect 5160 5646 5362 5650
rect 5436 5643 5444 5650
rect 5550 5643 5558 5821
rect 5872 5786 5885 5838
rect 5937 5786 5950 5838
rect 5872 5774 5950 5786
rect 5872 5722 5885 5774
rect 5937 5722 5950 5774
rect 5872 5710 5950 5722
rect 5872 5658 5885 5710
rect 5937 5658 5950 5710
rect 5436 5614 5558 5643
rect 5678 5638 5756 5650
rect 5678 5586 5691 5638
rect 5743 5586 5756 5638
rect 5678 5574 5756 5586
rect 5678 5522 5691 5574
rect 5743 5522 5756 5574
rect 5678 5510 5756 5522
rect 5872 5646 5950 5658
rect 5872 5594 5885 5646
rect 5937 5594 5950 5646
rect 5872 5582 5950 5594
rect 5872 5530 5885 5582
rect 5937 5530 5950 5582
rect 5872 5520 5950 5530
rect 6064 5964 6142 5974
rect 6064 5912 6077 5964
rect 6129 5912 6142 5964
rect 6064 5900 6142 5912
rect 6064 5848 6077 5900
rect 6129 5848 6142 5900
rect 6064 5836 6142 5848
rect 6064 5784 6077 5836
rect 6129 5784 6142 5836
rect 6064 5772 6142 5784
rect 6064 5720 6077 5772
rect 6129 5720 6142 5772
rect 6064 5708 6142 5720
rect 6064 5656 6077 5708
rect 6129 5656 6142 5708
rect 6064 5644 6142 5656
rect 6064 5592 6077 5644
rect 6129 5592 6142 5644
rect 6064 5580 6142 5592
rect 6064 5528 6077 5580
rect 6129 5528 6142 5580
rect 6064 5518 6142 5528
rect 6256 5950 6334 5960
rect 6256 5898 6269 5950
rect 6321 5898 6334 5950
rect 6256 5886 6334 5898
rect 6256 5834 6269 5886
rect 6321 5834 6334 5886
rect 6256 5822 6334 5834
rect 6256 5770 6269 5822
rect 6321 5770 6334 5822
rect 6256 5758 6334 5770
rect 6256 5706 6269 5758
rect 6321 5706 6334 5758
rect 6256 5694 6334 5706
rect 6256 5642 6269 5694
rect 6321 5642 6334 5694
rect 6256 5630 6334 5642
rect 6256 5578 6269 5630
rect 6321 5578 6334 5630
rect 6256 5566 6334 5578
rect 6256 5514 6269 5566
rect 6321 5514 6334 5566
rect 6256 5504 6334 5514
rect 6448 5950 6526 5960
rect 6448 5898 6461 5950
rect 6513 5898 6526 5950
rect 6448 5886 6526 5898
rect 6448 5834 6461 5886
rect 6513 5834 6526 5886
rect 6448 5822 6526 5834
rect 6448 5770 6461 5822
rect 6513 5770 6526 5822
rect 6448 5758 6526 5770
rect 6448 5706 6461 5758
rect 6513 5706 6526 5758
rect 6448 5694 6526 5706
rect 6448 5642 6461 5694
rect 6513 5642 6526 5694
rect 6448 5630 6526 5642
rect 6448 5578 6461 5630
rect 6513 5578 6526 5630
rect 6448 5566 6526 5578
rect 6448 5514 6461 5566
rect 6513 5514 6526 5566
rect 6448 5504 6526 5514
rect 6886 5454 6968 7112
rect 7564 7088 7575 7268
rect 7755 7160 7818 7268
rect 7755 7088 7816 7160
rect 8882 7144 8966 7148
rect 7564 6914 7816 7088
rect 8048 7113 8162 7134
rect 8048 7061 8079 7113
rect 8131 7061 8162 7113
rect 8048 7049 8162 7061
rect 8048 6997 8079 7049
rect 8131 6997 8162 7049
rect 8504 7113 8580 7140
rect 8504 7061 8516 7113
rect 8568 7061 8580 7113
rect 8504 7034 8580 7061
rect 8692 7115 8768 7142
rect 8692 7063 8704 7115
rect 8756 7063 8768 7115
rect 8692 7036 8768 7063
rect 8882 7092 8898 7144
rect 8950 7092 8966 7144
rect 8882 7080 8966 7092
rect 8882 7028 8898 7080
rect 8950 7028 8966 7080
rect 8882 7024 8966 7028
rect 8048 6976 8162 6997
rect 9002 6962 9092 7420
rect 9236 7346 9528 7724
rect 9234 7321 9528 7346
rect 9234 7269 9281 7321
rect 9333 7269 9345 7321
rect 9397 7269 9528 7321
rect 10862 7310 10980 7326
rect 9234 7200 9528 7269
rect 9236 7190 9528 7200
rect 9950 7257 10054 7276
rect 9950 7205 9976 7257
rect 10028 7205 10054 7257
rect 10862 7258 10895 7310
rect 10947 7258 10980 7310
rect 10862 7242 10980 7258
rect 9240 7180 9436 7190
rect 9950 7186 10054 7205
rect 7558 6910 7956 6914
rect 7558 6906 8238 6910
rect 8372 6906 9092 6962
rect 9244 6978 9436 7180
rect 11630 7156 11830 7290
rect 11268 7146 11832 7156
rect 11268 7112 11291 7146
rect 11325 7112 11832 7146
rect 11268 7108 11832 7112
rect 11268 7102 11348 7108
rect 10912 7098 10960 7100
rect 10900 7090 10980 7098
rect 11630 7092 11830 7108
rect 10900 7038 10914 7090
rect 10966 7038 10980 7090
rect 10900 7030 10980 7038
rect 10122 7018 10350 7022
rect 10110 7012 10350 7018
rect 10110 6978 10122 7012
rect 10156 6996 10350 7012
rect 11072 7017 11158 7030
rect 11072 6996 11098 7017
rect 10156 6984 11098 6996
rect 10156 6978 10228 6984
rect 9244 6958 9494 6978
rect 10110 6972 10228 6978
rect 10296 6983 11098 6984
rect 11132 6983 11158 7017
rect 10296 6970 11158 6983
rect 10296 6968 11150 6970
rect 9244 6950 9896 6958
rect 9244 6941 10078 6950
rect 9244 6912 10021 6941
rect 7558 6902 9092 6906
rect 9216 6907 10021 6912
rect 10055 6907 10078 6941
rect 7558 6898 9088 6902
rect 7558 6850 8438 6898
rect 8766 6896 8980 6898
rect 9216 6896 10078 6907
rect 7558 6840 8404 6850
rect 9216 6842 9896 6896
rect 7558 6838 8238 6840
rect 7840 6834 8238 6838
rect 7960 6779 8124 6792
rect 7960 6727 7984 6779
rect 8036 6727 8048 6779
rect 8100 6727 8124 6779
rect 9216 6748 9522 6842
rect 10856 6772 11006 6790
rect 10824 6764 11006 6772
rect 7960 6714 8124 6727
rect 9012 6662 9552 6748
rect 9010 6580 9552 6662
rect 9938 6718 10070 6760
rect 10824 6724 10873 6764
rect 9938 6666 9972 6718
rect 10024 6666 10070 6718
rect 10856 6712 10873 6724
rect 10925 6712 10937 6764
rect 10989 6712 11006 6764
rect 10856 6686 11006 6712
rect 9938 6660 10070 6666
rect 9952 6640 9962 6660
rect 7344 6502 8634 6504
rect 9010 6502 9092 6580
rect 9428 6566 9500 6580
rect 10334 6540 10492 6548
rect 10334 6524 10355 6540
rect 7344 6420 9092 6502
rect 10332 6488 10355 6524
rect 10407 6488 10419 6540
rect 10471 6524 10492 6540
rect 10471 6488 10496 6524
rect 10332 6482 10361 6488
rect 10395 6482 10433 6488
rect 10467 6482 10496 6488
rect 10332 6474 10496 6482
rect 10434 6434 12558 6444
rect 7344 6418 9034 6420
rect 7344 6416 8634 6418
rect 7346 6350 7454 6416
rect 8278 6377 8352 6382
rect 7346 6302 7782 6350
rect 7348 6284 7782 6302
rect 8278 6325 8289 6377
rect 8341 6325 8352 6377
rect 8278 6313 8352 6325
rect 7348 6026 7452 6284
rect 8278 6261 8289 6313
rect 8341 6261 8352 6313
rect 8278 6256 8352 6261
rect 8470 6377 8544 6382
rect 8470 6325 8481 6377
rect 8533 6325 8544 6377
rect 9634 6362 12558 6434
rect 9634 6358 9714 6362
rect 8470 6313 8544 6325
rect 8470 6261 8481 6313
rect 8533 6261 8544 6313
rect 8674 6344 8770 6354
rect 8674 6292 8696 6344
rect 8748 6292 8770 6344
rect 8674 6282 8770 6292
rect 9586 6332 9714 6358
rect 8470 6256 8544 6261
rect 7784 6226 7870 6234
rect 7784 6174 7801 6226
rect 7853 6174 7870 6226
rect 9586 6176 9698 6332
rect 9580 6174 9728 6176
rect 7784 6166 7870 6174
rect 8958 6170 9728 6174
rect 7502 6122 7588 6142
rect 7502 6070 7519 6122
rect 7571 6070 7588 6122
rect 7502 6058 7588 6070
rect 8168 6122 8254 6142
rect 8168 6070 8185 6122
rect 8237 6070 8254 6122
rect 8168 6058 8254 6070
rect 8366 6120 8452 6140
rect 8366 6068 8383 6120
rect 8435 6068 8452 6120
rect 8366 6056 8452 6068
rect 8562 6138 8648 6142
rect 8948 6138 9728 6170
rect 8562 6122 9728 6138
rect 10584 6136 10688 6140
rect 8562 6070 8579 6122
rect 8631 6098 9728 6122
rect 8631 6094 9414 6098
rect 8631 6070 9042 6094
rect 8562 6058 9042 6070
rect 8578 6046 9042 6058
rect 9368 6057 9454 6062
rect 8948 6028 9040 6046
rect 7348 6002 7458 6026
rect 7348 5946 7798 6002
rect 7350 5944 7798 5946
rect 7350 5758 7458 5944
rect 8960 5838 9024 6028
rect 9368 6005 9385 6057
rect 9437 6005 9454 6057
rect 9368 6000 9454 6005
rect 9580 5960 9728 6098
rect 9104 5926 9176 5932
rect 9104 5874 9114 5926
rect 9166 5874 9176 5926
rect 9582 5892 9728 5960
rect 9104 5868 9176 5874
rect 8944 5758 9400 5838
rect 7350 5664 8738 5758
rect 9016 5726 9218 5730
rect 9014 5720 9218 5726
rect 9014 5709 9055 5720
rect 9107 5709 9119 5720
rect 9171 5709 9218 5720
rect 9014 5675 9028 5709
rect 9171 5675 9172 5709
rect 9206 5675 9218 5709
rect 9014 5668 9055 5675
rect 9107 5668 9119 5675
rect 9171 5668 9218 5675
rect 7350 5654 7458 5664
rect 9014 5662 9218 5668
rect 9016 5654 9218 5662
rect 5626 5448 6276 5454
rect 6358 5448 6968 5454
rect 5626 5380 6968 5448
rect 6254 5192 6336 5380
rect 6366 5370 6968 5380
rect 7874 5385 8132 5398
rect 7874 5205 7923 5385
rect 8103 5205 8132 5385
rect 7874 5192 8132 5205
rect 4222 5100 4316 5124
rect 4014 5048 4243 5100
rect 4295 5048 4360 5100
rect 4014 5016 4360 5048
rect 4598 5088 6338 5192
rect 4598 4790 4678 5088
rect 6254 4968 6336 5088
rect 5964 4916 6336 4968
rect 5964 4900 6356 4916
rect 6136 4860 6214 4862
rect 6024 4858 6102 4860
rect 6024 4806 6037 4858
rect 6089 4806 6102 4858
rect 6136 4808 6149 4860
rect 6201 4808 6214 4860
rect 6136 4806 6214 4808
rect 6024 4804 6102 4806
rect 3566 4774 4354 4788
rect 4430 4786 4680 4790
rect 3566 4740 4292 4774
rect 4326 4740 4354 4774
rect 3566 4712 4354 4740
rect 4418 4777 4680 4786
rect 4418 4743 4441 4777
rect 4475 4774 4680 4777
rect 4475 4743 4682 4774
rect 4418 4734 4682 4743
rect 4434 4730 4682 4734
rect 5916 4738 5994 4740
rect 5916 4686 5929 4738
rect 5981 4686 5994 4738
rect 5916 4684 5994 4686
rect 6274 4642 6356 4900
rect 9580 4700 9728 5892
rect 10062 6074 10091 6126
rect 10143 6074 10172 6126
rect 10062 6062 10172 6074
rect 10062 6010 10091 6062
rect 10143 6010 10172 6062
rect 10062 5998 10172 6010
rect 10062 5946 10091 5998
rect 10143 5946 10172 5998
rect 10062 5934 10172 5946
rect 10062 5882 10091 5934
rect 10143 5882 10172 5934
rect 10398 5876 10408 6120
rect 10584 6084 10610 6136
rect 10662 6084 10688 6136
rect 11100 6120 11204 6124
rect 10584 6072 10688 6084
rect 10584 6020 10610 6072
rect 10662 6020 10688 6072
rect 10584 6008 10688 6020
rect 10584 5956 10610 6008
rect 10662 5956 10688 6008
rect 10584 5944 10688 5956
rect 10584 5892 10610 5944
rect 10662 5892 10688 5944
rect 10584 5888 10688 5892
rect 10914 5876 10924 6120
rect 11100 6068 11126 6120
rect 11178 6068 11204 6120
rect 11100 6056 11204 6068
rect 11100 6004 11126 6056
rect 11178 6004 11204 6056
rect 11100 5992 11204 6004
rect 11100 5940 11126 5992
rect 11178 5940 11204 5992
rect 11100 5928 11204 5940
rect 11100 5876 11126 5928
rect 11178 5876 11204 5928
rect 11428 5890 11438 6134
rect 12642 6126 12746 6130
rect 11618 6112 11722 6116
rect 12130 6112 12234 6116
rect 11618 6060 11644 6112
rect 11696 6060 11722 6112
rect 11618 6048 11722 6060
rect 11618 5996 11644 6048
rect 11696 5996 11722 6048
rect 11618 5984 11722 5996
rect 11618 5932 11644 5984
rect 11696 5932 11722 5984
rect 11618 5920 11722 5932
rect 11100 5872 11204 5876
rect 11618 5868 11644 5920
rect 11696 5868 11722 5920
rect 11944 5868 11954 6112
rect 12130 6060 12156 6112
rect 12208 6060 12234 6112
rect 12130 6048 12234 6060
rect 12130 5996 12156 6048
rect 12208 5996 12234 6048
rect 12130 5984 12234 5996
rect 12130 5932 12156 5984
rect 12208 5932 12234 5984
rect 12130 5920 12234 5932
rect 12130 5868 12156 5920
rect 12208 5868 12234 5920
rect 12642 6074 12668 6126
rect 12720 6074 12746 6126
rect 12642 6062 12746 6074
rect 12642 6010 12668 6062
rect 12720 6010 12746 6062
rect 12642 5998 12746 6010
rect 12642 5946 12668 5998
rect 12720 5946 12746 5998
rect 12642 5934 12746 5946
rect 12642 5882 12668 5934
rect 12720 5882 12746 5934
rect 12642 5878 12746 5882
rect 11618 5864 11722 5868
rect 12130 5864 12234 5868
rect 10332 5122 10408 5188
rect 10836 5127 10960 5142
rect 10330 5113 10426 5122
rect 10330 5061 10352 5113
rect 10404 5061 10426 5113
rect 10330 5049 10426 5061
rect 10330 4997 10352 5049
rect 10404 4997 10426 5049
rect 10330 4985 10426 4997
rect 10330 4933 10352 4985
rect 10404 4933 10426 4985
rect 10330 4924 10426 4933
rect 10836 5075 10872 5127
rect 10924 5075 10960 5127
rect 10836 5063 10960 5075
rect 10836 5011 10872 5063
rect 10924 5011 10960 5063
rect 10836 4999 10960 5011
rect 10836 4947 10872 4999
rect 10924 4947 10960 4999
rect 10836 4932 10960 4947
rect 11360 5113 11484 5128
rect 11360 5061 11396 5113
rect 11448 5061 11484 5113
rect 11360 5049 11484 5061
rect 11360 4997 11396 5049
rect 11448 4997 11484 5049
rect 11360 4985 11484 4997
rect 11360 4933 11396 4985
rect 11448 4933 11484 4985
rect 11360 4918 11484 4933
rect 11864 5123 11988 5138
rect 11864 5071 11900 5123
rect 11952 5071 11988 5123
rect 11864 5059 11988 5071
rect 11864 5007 11900 5059
rect 11952 5007 11988 5059
rect 11864 4995 11988 5007
rect 11864 4943 11900 4995
rect 11952 4943 11988 4995
rect 11864 4928 11988 4943
rect 12382 5127 12506 5142
rect 12382 5075 12418 5127
rect 12470 5075 12506 5127
rect 12382 5063 12506 5075
rect 12382 5011 12418 5063
rect 12470 5011 12506 5063
rect 12382 4999 12506 5011
rect 12382 4947 12418 4999
rect 12470 4947 12506 4999
rect 12382 4932 12506 4947
rect 5944 4560 6356 4642
rect 9544 4616 12570 4700
rect 4070 4539 4314 4556
rect 4070 4487 4241 4539
rect 4293 4487 4314 4539
rect 4070 4476 4314 4487
rect 4220 4474 4314 4476
<< via1 >>
rect 6800 10739 6980 10919
rect 10711 11656 10763 11708
rect 10775 11656 10827 11708
rect 10839 11656 10891 11708
rect 10903 11656 10955 11708
rect 10967 11656 11019 11708
rect 11031 11656 11083 11708
rect 11095 11656 11147 11708
rect 11159 11656 11211 11708
rect 11223 11656 11275 11708
rect 11287 11656 11339 11708
rect 11351 11656 11403 11708
rect 11415 11656 11467 11708
rect 11479 11656 11531 11708
rect 11744 11555 11796 11607
rect 11808 11555 11860 11607
rect 11872 11555 11924 11607
rect 11936 11555 11988 11607
rect 12000 11555 12052 11607
rect 12064 11555 12116 11607
rect 12128 11555 12180 11607
rect 10715 11462 10767 11514
rect 10779 11462 10831 11514
rect 10843 11462 10895 11514
rect 10907 11462 10959 11514
rect 10971 11462 11023 11514
rect 11035 11462 11087 11514
rect 11099 11462 11151 11514
rect 11163 11462 11215 11514
rect 11227 11462 11279 11514
rect 11291 11462 11343 11514
rect 11355 11462 11407 11514
rect 11419 11462 11471 11514
rect 11483 11462 11535 11514
rect 11736 11367 11788 11419
rect 11800 11367 11852 11419
rect 11864 11367 11916 11419
rect 11928 11367 11980 11419
rect 11992 11367 12044 11419
rect 12056 11367 12108 11419
rect 12120 11367 12172 11419
rect 10725 11262 10777 11314
rect 10789 11262 10841 11314
rect 10853 11262 10905 11314
rect 10917 11262 10969 11314
rect 10981 11262 11033 11314
rect 11045 11262 11097 11314
rect 11109 11262 11161 11314
rect 11173 11262 11225 11314
rect 11237 11262 11289 11314
rect 11301 11262 11353 11314
rect 11365 11262 11417 11314
rect 11429 11262 11481 11314
rect 11493 11262 11545 11314
rect 11853 11176 12097 11177
rect 11853 10998 12097 11176
rect 11853 10997 12097 10998
rect 4847 9953 5091 10325
rect 5499 10313 5551 10365
rect 5499 10249 5551 10301
rect 5499 10185 5551 10237
rect 5499 10121 5551 10173
rect 5499 10057 5551 10109
rect 5499 9993 5551 10045
rect 6561 10315 6613 10367
rect 6561 10251 6613 10303
rect 6561 10187 6613 10239
rect 6561 10123 6613 10175
rect 6676 10197 6728 10249
rect 6676 10133 6728 10185
rect 6561 10059 6613 10111
rect 6561 9995 6613 10047
rect 7586 9952 7638 10004
rect 7586 9888 7638 9940
rect 7788 9950 7840 10002
rect 7788 9886 7840 9938
rect 7976 9956 8028 10008
rect 7976 9892 8028 9944
rect 4843 9315 5087 9687
rect 5517 9161 5569 9213
rect 5517 9097 5569 9149
rect 5517 9033 5569 9085
rect 6581 9127 6633 9179
rect 6581 9063 6633 9115
rect 6703 9104 6755 9156
rect 6581 8999 6633 9051
rect 6703 9040 6755 9092
rect 7686 8918 7738 8970
rect 7686 8854 7738 8906
rect 7884 8912 7936 8964
rect 7884 8848 7936 8900
rect 8100 8929 8152 8945
rect 8100 8895 8106 8929
rect 8106 8895 8140 8929
rect 8140 8895 8152 8929
rect 8100 8893 8152 8895
rect 5543 8109 5595 8161
rect 5543 8045 5595 8097
rect 5543 7981 5595 8033
rect 5543 7917 5595 7969
rect 5543 7853 5595 7905
rect 6606 8046 6658 8098
rect 6606 7982 6658 8034
rect 6730 7994 6782 8046
rect 6606 7918 6658 7970
rect 6730 7930 6782 7982
rect 5543 7789 5595 7841
rect 4371 7539 4551 7719
rect 7887 8251 7896 8258
rect 7896 8251 7930 8258
rect 7930 8251 7939 8258
rect 7887 8213 7939 8251
rect 7887 8206 7896 8213
rect 7896 8206 7930 8213
rect 7930 8206 7939 8213
rect 9249 10308 9621 10488
rect 9749 9594 9801 9646
rect 9947 9588 9999 9640
rect 10133 9586 10185 9638
rect 10364 9614 10416 9636
rect 10364 9584 10398 9614
rect 10398 9584 10416 9614
rect 11628 9469 11872 9841
rect 9849 9358 9901 9410
rect 10039 9356 10091 9408
rect 10231 9360 10283 9412
rect 11625 8829 11869 9201
rect 8358 8147 8410 8199
rect 8422 8147 8474 8199
rect 9221 7905 9273 7957
rect 9221 7841 9273 7893
rect 9221 7777 9273 7829
rect 14286 7909 14338 7961
rect 14286 7845 14338 7897
rect 14286 7781 14338 7833
rect 4642 6755 4886 7127
rect 4642 6085 4886 6457
rect 7947 7365 7999 7417
rect 7947 7301 7999 7353
rect 8410 7299 8462 7351
rect 8602 7297 8654 7349
rect 8804 7295 8856 7347
rect 5595 7018 5647 7070
rect 5595 6954 5647 7006
rect 5595 6890 5647 6942
rect 5595 6826 5647 6878
rect 5595 6762 5647 6814
rect 5595 6698 5647 6750
rect 5595 6634 5647 6686
rect 5787 7014 5839 7066
rect 5787 6950 5839 7002
rect 5787 6886 5839 6938
rect 5787 6822 5839 6874
rect 5787 6758 5839 6810
rect 5787 6694 5839 6746
rect 5787 6630 5839 6682
rect 5981 7020 6033 7072
rect 5981 6956 6033 7008
rect 5981 6892 6033 6944
rect 5981 6828 6033 6880
rect 5981 6764 6033 6816
rect 5981 6700 6033 6752
rect 5981 6636 6033 6688
rect 6173 7018 6225 7070
rect 6173 6954 6225 7006
rect 6173 6890 6225 6942
rect 6173 6826 6225 6878
rect 6173 6762 6225 6814
rect 6173 6698 6225 6750
rect 6173 6634 6225 6686
rect 6367 7018 6419 7070
rect 6367 6954 6419 7006
rect 6367 6890 6419 6942
rect 6367 6826 6419 6878
rect 6367 6762 6419 6814
rect 6367 6698 6419 6750
rect 6367 6634 6419 6686
rect 6559 7014 6611 7066
rect 6559 6950 6611 7002
rect 6559 6886 6611 6938
rect 6559 6822 6611 6874
rect 6559 6758 6611 6810
rect 6559 6694 6611 6746
rect 6559 6630 6611 6682
rect 5691 5910 5743 5962
rect 5691 5846 5743 5898
rect 5885 5914 5937 5966
rect 5885 5850 5937 5902
rect 5473 5821 5525 5832
rect 5473 5780 5525 5821
rect 5473 5716 5525 5768
rect 5473 5652 5525 5704
rect 5885 5786 5937 5838
rect 5885 5722 5937 5774
rect 5885 5658 5937 5710
rect 5691 5586 5743 5638
rect 5691 5522 5743 5574
rect 5885 5594 5937 5646
rect 5885 5530 5937 5582
rect 6077 5912 6129 5964
rect 6077 5848 6129 5900
rect 6077 5784 6129 5836
rect 6077 5720 6129 5772
rect 6077 5656 6129 5708
rect 6077 5592 6129 5644
rect 6077 5528 6129 5580
rect 6269 5898 6321 5950
rect 6269 5834 6321 5886
rect 6269 5770 6321 5822
rect 6269 5706 6321 5758
rect 6269 5642 6321 5694
rect 6269 5578 6321 5630
rect 6269 5514 6321 5566
rect 6461 5898 6513 5950
rect 6461 5834 6513 5886
rect 6461 5770 6513 5822
rect 6461 5706 6513 5758
rect 6461 5642 6513 5694
rect 6461 5578 6513 5630
rect 6461 5514 6513 5566
rect 7575 7088 7755 7268
rect 8079 7061 8131 7113
rect 8079 6997 8131 7049
rect 8516 7061 8568 7113
rect 8704 7063 8756 7115
rect 8898 7092 8950 7144
rect 8898 7028 8950 7080
rect 9281 7269 9333 7321
rect 9345 7269 9397 7321
rect 9976 7205 10028 7257
rect 10895 7258 10947 7310
rect 10914 7086 10966 7090
rect 10914 7052 10919 7086
rect 10919 7052 10953 7086
rect 10953 7052 10966 7086
rect 10914 7038 10966 7052
rect 7984 6727 8036 6779
rect 8048 6727 8100 6779
rect 9972 6666 10024 6718
rect 10873 6712 10925 6764
rect 10937 6712 10989 6764
rect 10355 6516 10407 6540
rect 10355 6488 10361 6516
rect 10361 6488 10395 6516
rect 10395 6488 10407 6516
rect 10419 6516 10471 6540
rect 10419 6488 10433 6516
rect 10433 6488 10467 6516
rect 10467 6488 10471 6516
rect 8289 6325 8341 6377
rect 8289 6261 8341 6313
rect 8481 6325 8533 6377
rect 8481 6261 8533 6313
rect 8696 6292 8748 6344
rect 7801 6174 7853 6226
rect 7519 6070 7571 6122
rect 8185 6070 8237 6122
rect 8383 6068 8435 6120
rect 8579 6070 8631 6122
rect 9385 6005 9437 6057
rect 9114 5874 9166 5926
rect 9055 5709 9107 5720
rect 9119 5709 9171 5720
rect 9055 5675 9062 5709
rect 9062 5675 9100 5709
rect 9100 5675 9107 5709
rect 9119 5675 9134 5709
rect 9134 5675 9171 5709
rect 9055 5668 9107 5675
rect 9119 5668 9171 5675
rect 7923 5205 8103 5385
rect 4243 5048 4295 5100
rect 6037 4806 6089 4858
rect 6149 4808 6201 4860
rect 5929 4686 5981 4738
rect 10091 6074 10143 6126
rect 10091 6010 10143 6062
rect 10091 5946 10143 5998
rect 10091 5882 10143 5934
rect 10610 6084 10662 6136
rect 10610 6020 10662 6072
rect 10610 5956 10662 6008
rect 10610 5892 10662 5944
rect 11126 6068 11178 6120
rect 11126 6004 11178 6056
rect 11126 5940 11178 5992
rect 11126 5876 11178 5928
rect 11644 6060 11696 6112
rect 11644 5996 11696 6048
rect 11644 5932 11696 5984
rect 11644 5868 11696 5920
rect 12156 6060 12208 6112
rect 12156 5996 12208 6048
rect 12156 5932 12208 5984
rect 12156 5868 12208 5920
rect 12668 6074 12720 6126
rect 12668 6010 12720 6062
rect 12668 5946 12720 5998
rect 12668 5882 12720 5934
rect 10352 5061 10404 5113
rect 10352 4997 10404 5049
rect 10352 4933 10404 4985
rect 10872 5075 10924 5127
rect 10872 5011 10924 5063
rect 10872 4947 10924 4999
rect 11396 5061 11448 5113
rect 11396 4997 11448 5049
rect 11396 4933 11448 4985
rect 11900 5071 11952 5123
rect 11900 5007 11952 5059
rect 11900 4943 11952 4995
rect 12418 5075 12470 5127
rect 12418 5011 12470 5063
rect 12418 4947 12470 4999
rect 4241 4487 4293 4539
<< metal2 >>
rect 10694 11708 11548 11718
rect 10694 11656 10711 11708
rect 10763 11656 10775 11708
rect 10827 11656 10839 11708
rect 10891 11656 10903 11708
rect 10955 11656 10967 11708
rect 11019 11656 11031 11708
rect 11083 11656 11095 11708
rect 11147 11656 11159 11708
rect 11211 11656 11223 11708
rect 11275 11656 11287 11708
rect 11339 11656 11351 11708
rect 11403 11656 11415 11708
rect 11467 11656 11479 11708
rect 11531 11656 11548 11708
rect 10694 11646 11548 11656
rect 10928 11524 11258 11646
rect 11734 11607 12190 11618
rect 11734 11555 11744 11607
rect 11796 11555 11808 11607
rect 11860 11555 11872 11607
rect 11924 11555 11936 11607
rect 11988 11555 12000 11607
rect 12052 11555 12064 11607
rect 12116 11555 12128 11607
rect 12180 11555 12190 11607
rect 11734 11544 12190 11555
rect 10698 11514 11552 11524
rect 10698 11462 10715 11514
rect 10767 11462 10779 11514
rect 10831 11462 10843 11514
rect 10895 11462 10907 11514
rect 10959 11462 10971 11514
rect 11023 11462 11035 11514
rect 11087 11462 11099 11514
rect 11151 11462 11163 11514
rect 11215 11462 11227 11514
rect 11279 11462 11291 11514
rect 11343 11462 11355 11514
rect 11407 11462 11419 11514
rect 11471 11462 11483 11514
rect 11535 11462 11552 11514
rect 10698 11452 11552 11462
rect 10928 11324 11258 11452
rect 11846 11430 12104 11544
rect 11726 11419 12182 11430
rect 11726 11367 11736 11419
rect 11788 11367 11800 11419
rect 11852 11367 11864 11419
rect 11916 11367 11928 11419
rect 11980 11367 11992 11419
rect 12044 11367 12056 11419
rect 12108 11367 12120 11419
rect 12172 11367 12182 11419
rect 11726 11356 12182 11367
rect 10708 11314 11562 11324
rect 10708 11262 10725 11314
rect 10777 11262 10789 11314
rect 10841 11262 10853 11314
rect 10905 11262 10917 11314
rect 10969 11262 10981 11314
rect 11033 11262 11045 11314
rect 11097 11262 11109 11314
rect 11161 11262 11173 11314
rect 11225 11262 11237 11314
rect 11289 11262 11301 11314
rect 11353 11262 11365 11314
rect 11417 11262 11429 11314
rect 11481 11262 11493 11314
rect 11545 11262 11562 11314
rect 10708 11252 11562 11262
rect 10928 11118 11258 11252
rect 11846 11206 12104 11356
rect 11840 11177 12110 11206
rect 6782 10919 6998 10946
rect 6782 10897 6800 10919
rect 6980 10918 6998 10919
rect 6980 10897 7008 10918
rect 6998 10761 7008 10897
rect 6782 10739 6800 10761
rect 6980 10739 7008 10761
rect 6782 10710 7008 10739
rect 10959 10538 11197 11118
rect 11840 10997 11853 11177
rect 12097 10997 12110 11177
rect 11840 10968 12110 10997
rect 11846 10958 12104 10968
rect 9242 10512 9628 10516
rect 10928 10512 11258 10538
rect 8434 10488 11264 10512
rect 5494 10365 5556 10388
rect 4840 10325 5098 10356
rect 4840 9953 4847 10325
rect 5091 9953 5098 10325
rect 5494 10313 5499 10365
rect 5551 10313 5556 10365
rect 5494 10301 5556 10313
rect 5494 10249 5499 10301
rect 5551 10249 5556 10301
rect 6560 10367 6614 10388
rect 6560 10315 6561 10367
rect 6613 10315 6614 10367
rect 6560 10303 6614 10315
rect 6560 10300 6561 10303
rect 5494 10237 5556 10249
rect 5494 10185 5499 10237
rect 5551 10185 5556 10237
rect 5494 10173 5556 10185
rect 5494 10121 5499 10173
rect 5551 10121 5556 10173
rect 5494 10109 5556 10121
rect 6558 10251 6561 10300
rect 6613 10300 6614 10303
rect 8434 10308 9249 10488
rect 9621 10308 11264 10488
rect 8434 10300 11264 10308
rect 6613 10276 6628 10300
rect 6558 10239 6565 10251
rect 6558 10187 6561 10239
rect 6621 10220 6628 10276
rect 6682 10272 6752 10292
rect 6613 10196 6628 10220
rect 6558 10175 6565 10187
rect 6558 10123 6561 10175
rect 6621 10140 6628 10196
rect 6613 10123 6628 10140
rect 6558 10116 6628 10123
rect 6672 10268 6752 10272
rect 6672 10249 6689 10268
rect 6672 10197 6676 10249
rect 6745 10212 6752 10268
rect 6728 10197 6752 10212
rect 6672 10188 6752 10197
rect 6672 10185 6689 10188
rect 6672 10133 6676 10185
rect 6672 10132 6689 10133
rect 6745 10132 6752 10188
rect 5494 10057 5499 10109
rect 5551 10057 5556 10109
rect 5494 10045 5556 10057
rect 5494 9993 5499 10045
rect 5551 9993 5556 10045
rect 5494 9970 5556 9993
rect 6560 10111 6614 10116
rect 6560 10059 6561 10111
rect 6613 10059 6614 10111
rect 6672 10110 6752 10132
rect 6682 10108 6752 10110
rect 8434 10084 8646 10300
rect 9242 10280 9628 10300
rect 6560 10047 6614 10059
rect 6560 9995 6561 10047
rect 6613 9995 6614 10047
rect 7596 10034 8646 10084
rect 6560 9974 6614 9995
rect 7586 10008 8646 10034
rect 7586 10004 7976 10008
rect 4840 9944 4869 9953
rect 5085 9944 5098 9953
rect 4840 9922 5098 9944
rect 7638 10002 7976 10004
rect 7638 9952 7788 10002
rect 7586 9950 7788 9952
rect 7840 9956 7976 10002
rect 8028 9956 8646 10008
rect 7840 9950 8646 9956
rect 7586 9944 8646 9950
rect 7586 9940 7976 9944
rect 7638 9938 7976 9940
rect 7638 9888 7788 9938
rect 7586 9886 7788 9888
rect 7840 9892 7976 9938
rect 8028 9892 8646 9944
rect 7840 9886 8646 9892
rect 7586 9872 8646 9886
rect 7586 9858 7638 9872
rect 7788 9856 7840 9872
rect 7976 9862 8028 9872
rect 11622 9849 11874 9878
rect 11622 9841 11640 9849
rect 11856 9841 11874 9849
rect 4836 9687 5094 9718
rect 4836 9315 4843 9687
rect 5087 9315 5094 9687
rect 4836 9284 5094 9315
rect 9712 9682 9786 9702
rect 9712 9676 9812 9682
rect 9712 9646 10196 9676
rect 9712 9594 9749 9646
rect 9801 9640 10196 9646
rect 9801 9594 9947 9640
rect 9712 9588 9947 9594
rect 9999 9638 10196 9640
rect 9999 9588 10133 9638
rect 9712 9586 10133 9588
rect 10185 9586 10196 9638
rect 9712 9568 10196 9586
rect 10356 9638 10424 9670
rect 10356 9582 10362 9638
rect 10418 9582 10424 9638
rect 9712 9558 9812 9568
rect 5516 9213 5570 9254
rect 5516 9161 5517 9213
rect 5569 9161 5570 9213
rect 5516 9149 5570 9161
rect 5516 9097 5517 9149
rect 5569 9097 5570 9149
rect 5516 9085 5570 9097
rect 5516 9033 5517 9085
rect 5569 9033 5570 9085
rect 5516 8992 5570 9033
rect 6568 9179 6646 9190
rect 6568 9127 6581 9179
rect 6633 9127 6646 9179
rect 6568 9115 6646 9127
rect 6568 9063 6581 9115
rect 6633 9063 6646 9115
rect 6568 9051 6646 9063
rect 6568 8999 6581 9051
rect 6633 8999 6646 9051
rect 6700 9156 6758 9182
rect 6700 9104 6703 9156
rect 6755 9104 6758 9156
rect 6700 9092 6758 9104
rect 6700 9040 6703 9092
rect 6755 9040 6758 9092
rect 6700 9014 6758 9040
rect 6568 8988 6646 8999
rect 7686 8988 7738 9000
rect 8096 8999 8172 9012
rect 7884 8988 7936 8994
rect 7686 8986 7940 8988
rect 8096 8986 8106 8999
rect 7686 8970 8106 8986
rect 7738 8964 8106 8970
rect 7738 8918 7884 8964
rect 7686 8912 7884 8918
rect 7936 8945 8106 8964
rect 8162 8986 8172 8999
rect 7936 8912 8100 8945
rect 8162 8943 8174 8986
rect 8152 8919 8174 8943
rect 7686 8906 8100 8912
rect 7738 8900 8100 8906
rect 7738 8854 7884 8900
rect 7686 8848 7884 8854
rect 7936 8893 8100 8900
rect 7936 8863 8106 8893
rect 8162 8863 8174 8919
rect 7936 8848 8174 8863
rect 7686 8836 8174 8848
rect 7686 8824 7738 8836
rect 7874 8834 8174 8836
rect 7884 8818 7936 8834
rect 9208 8478 9290 8488
rect 9712 8478 9786 9558
rect 9946 9552 10000 9568
rect 10132 9550 10186 9568
rect 10356 9550 10424 9582
rect 11622 9469 11628 9841
rect 11872 9469 11874 9841
rect 9838 9452 9912 9460
rect 9838 9415 10304 9452
rect 11622 9444 11874 9469
rect 11626 9434 11874 9444
rect 9838 9359 9847 9415
rect 9903 9412 10304 9415
rect 9903 9408 10231 9412
rect 9903 9359 10039 9408
rect 9838 9358 9849 9359
rect 9901 9358 10039 9359
rect 9838 9356 10039 9358
rect 10091 9360 10231 9408
rect 10283 9360 10304 9412
rect 10091 9356 10304 9360
rect 9838 9320 10304 9356
rect 9838 9314 9912 9320
rect 11606 9203 11888 9228
rect 11606 9201 11639 9203
rect 11855 9201 11888 9203
rect 11606 8829 11625 9201
rect 11869 8829 11888 9201
rect 11606 8827 11639 8829
rect 11855 8827 11888 8829
rect 11606 8802 11888 8827
rect 9198 8352 9852 8478
rect 7878 8260 7948 8296
rect 7878 8204 7885 8260
rect 7941 8204 7948 8260
rect 5538 8161 5600 8184
rect 7878 8168 7948 8204
rect 8348 8199 8484 8210
rect 5538 8109 5543 8161
rect 5595 8109 5600 8161
rect 8348 8147 8358 8199
rect 8410 8147 8422 8199
rect 8474 8147 8484 8199
rect 8348 8136 8484 8147
rect 5538 8097 5600 8109
rect 5538 8045 5543 8097
rect 5595 8045 5600 8097
rect 5538 8033 5600 8045
rect 5538 7981 5543 8033
rect 5595 7981 5600 8033
rect 5538 7969 5600 7981
rect 5538 7917 5543 7969
rect 5595 7917 5600 7969
rect 5538 7905 5600 7917
rect 5538 7853 5543 7905
rect 5595 7853 5600 7905
rect 6600 8098 6664 8128
rect 6600 8046 6606 8098
rect 6658 8046 6664 8098
rect 6600 8034 6664 8046
rect 6600 7982 6606 8034
rect 6658 7982 6664 8034
rect 6600 7970 6664 7982
rect 6600 7918 6606 7970
rect 6658 7918 6664 7970
rect 6600 7890 6664 7918
rect 6726 8046 6786 8062
rect 6726 7994 6730 8046
rect 6782 7994 6786 8046
rect 6726 7982 6786 7994
rect 6726 7930 6730 7982
rect 6782 7930 6786 7982
rect 9208 7964 9290 8352
rect 6726 7914 6786 7930
rect 7572 7957 9290 7964
rect 7572 7905 9221 7957
rect 9273 7905 9290 7957
rect 7572 7893 9290 7905
rect 6602 7880 6656 7890
rect 5538 7841 5600 7853
rect 5538 7789 5543 7841
rect 5595 7789 5600 7841
rect 5538 7766 5600 7789
rect 7572 7841 9221 7893
rect 9273 7841 9290 7893
rect 7572 7829 9290 7841
rect 7572 7777 9221 7829
rect 9273 7782 9290 7829
rect 14286 7961 14338 7974
rect 14338 7909 14352 7924
rect 14286 7897 14352 7909
rect 14338 7896 14352 7897
rect 14286 7840 14294 7845
rect 14350 7840 14352 7896
rect 14286 7833 14352 7840
rect 9273 7777 9286 7782
rect 7572 7756 9286 7777
rect 14338 7812 14352 7833
rect 14286 7768 14338 7781
rect 4364 7719 4558 7742
rect 4364 7539 4371 7719
rect 4551 7539 4558 7719
rect 4364 7516 4558 7539
rect 7580 7684 7766 7756
rect 9216 7752 9278 7756
rect 7074 7284 7196 7330
rect 7580 7298 7764 7684
rect 7926 7417 8020 7448
rect 7926 7392 7947 7417
rect 7574 7284 7764 7298
rect 7908 7365 7947 7392
rect 7999 7392 8020 7417
rect 7999 7384 8872 7392
rect 7999 7365 9442 7384
rect 7908 7353 9442 7365
rect 7908 7301 7947 7353
rect 7999 7351 9442 7353
rect 7999 7301 8410 7351
rect 7908 7299 8410 7301
rect 8462 7349 9442 7351
rect 8462 7299 8602 7349
rect 7908 7297 8602 7299
rect 8654 7347 9442 7349
rect 8654 7297 8804 7347
rect 7908 7295 8804 7297
rect 8856 7340 9442 7347
rect 8856 7321 9440 7340
rect 10876 7336 10990 7342
rect 8856 7295 9281 7321
rect 7908 7286 9281 7295
rect 7074 7268 7776 7284
rect 7926 7270 8020 7286
rect 4626 7127 4902 7168
rect 4626 6755 4642 7127
rect 4886 6755 4902 7127
rect 7074 7104 7575 7268
rect 5592 7070 5650 7090
rect 5592 7058 5595 7070
rect 4626 6714 4902 6755
rect 5562 7018 5595 7058
rect 5647 7058 5650 7070
rect 5784 7066 5842 7086
rect 5784 7058 5787 7066
rect 5647 7018 5787 7058
rect 5562 7014 5787 7018
rect 5839 7058 5842 7066
rect 5978 7072 6036 7092
rect 5978 7058 5981 7072
rect 5839 7020 5981 7058
rect 6033 7058 6036 7072
rect 6170 7070 6228 7090
rect 6170 7058 6173 7070
rect 6033 7020 6173 7058
rect 5839 7018 6173 7020
rect 6225 7058 6228 7070
rect 6364 7070 6422 7090
rect 6364 7058 6367 7070
rect 6225 7018 6367 7058
rect 6419 7058 6422 7070
rect 6556 7066 6614 7086
rect 6556 7058 6559 7066
rect 6419 7018 6559 7058
rect 5839 7014 6559 7018
rect 6611 7058 6614 7066
rect 6611 7014 6624 7058
rect 5562 7008 6624 7014
rect 5562 7006 5981 7008
rect 5562 6954 5595 7006
rect 5647 7002 5981 7006
rect 5647 6954 5787 7002
rect 5562 6950 5787 6954
rect 5839 6956 5981 7002
rect 6033 7006 6624 7008
rect 6033 6956 6173 7006
rect 5839 6954 6173 6956
rect 6225 6954 6367 7006
rect 6419 7002 6624 7006
rect 6419 6954 6559 7002
rect 5839 6950 6559 6954
rect 6611 6950 6624 7002
rect 5562 6944 6624 6950
rect 5562 6942 5981 6944
rect 5562 6890 5595 6942
rect 5647 6938 5981 6942
rect 5647 6890 5787 6938
rect 5562 6886 5787 6890
rect 5839 6892 5981 6938
rect 6033 6942 6624 6944
rect 6033 6892 6173 6942
rect 5839 6890 6173 6892
rect 6225 6890 6367 6942
rect 6419 6938 6624 6942
rect 6419 6890 6559 6938
rect 5839 6886 6559 6890
rect 6611 6886 6624 6938
rect 5562 6880 6624 6886
rect 5562 6878 5981 6880
rect 5562 6826 5595 6878
rect 5647 6874 5981 6878
rect 5647 6826 5787 6874
rect 5562 6822 5787 6826
rect 5839 6828 5981 6874
rect 6033 6878 6624 6880
rect 6033 6828 6173 6878
rect 5839 6826 6173 6828
rect 6225 6826 6367 6878
rect 6419 6874 6624 6878
rect 6419 6826 6559 6874
rect 5839 6822 6559 6826
rect 6611 6822 6624 6874
rect 5562 6816 6624 6822
rect 5562 6814 5981 6816
rect 5562 6762 5595 6814
rect 5647 6810 5981 6814
rect 5647 6762 5787 6810
rect 5562 6758 5787 6762
rect 5839 6764 5981 6810
rect 6033 6814 6624 6816
rect 7074 6844 7196 7104
rect 7574 7088 7575 7104
rect 7755 7104 7776 7268
rect 8408 7262 8464 7286
rect 8600 7260 8656 7286
rect 8802 7269 9281 7286
rect 9333 7269 9345 7321
rect 9397 7269 9440 7321
rect 10872 7313 10990 7336
rect 10872 7310 10905 7313
rect 8802 7264 9440 7269
rect 8802 7258 8858 7264
rect 9244 7208 9440 7264
rect 9960 7259 10044 7286
rect 9244 7180 9442 7208
rect 9960 7203 9974 7259
rect 10030 7203 10044 7259
rect 10872 7258 10895 7310
rect 10872 7257 10905 7258
rect 10961 7257 10990 7313
rect 10872 7232 10990 7257
rect 10876 7228 10990 7232
rect 9960 7176 10044 7203
rect 8892 7152 8956 7158
rect 8062 7144 8152 7148
rect 8058 7121 8152 7144
rect 7755 7094 7764 7104
rect 7755 7088 7756 7094
rect 7574 7064 7756 7088
rect 8058 7061 8079 7121
rect 8135 7065 8152 7121
rect 8131 7061 8152 7065
rect 8058 7049 8152 7061
rect 8058 6985 8079 7049
rect 8131 7041 8152 7049
rect 8135 6985 8152 7041
rect 8512 7144 8956 7152
rect 8512 7115 8898 7144
rect 8512 7113 8704 7115
rect 8512 7061 8516 7113
rect 8568 7063 8704 7113
rect 8756 7114 8898 7115
rect 8950 7114 8956 7144
rect 8756 7063 8896 7114
rect 8568 7061 8896 7063
rect 8512 7058 8896 7061
rect 8952 7070 8956 7114
rect 10910 7100 10970 7108
rect 10592 7090 10972 7100
rect 8952 7058 8964 7070
rect 8512 7028 8898 7058
rect 8950 7028 8964 7058
rect 10592 7038 10914 7090
rect 10966 7038 10972 7090
rect 10592 7028 10972 7038
rect 8514 7012 8574 7028
rect 8702 7026 8758 7028
rect 8892 7022 8962 7028
rect 8892 7014 8956 7022
rect 8058 6966 8152 6985
rect 8062 6958 8152 6966
rect 10594 6998 10676 7028
rect 10910 7020 10970 7028
rect 7074 6814 7194 6844
rect 6033 6764 6173 6814
rect 5839 6762 6173 6764
rect 6225 6762 6367 6814
rect 6419 6810 7196 6814
rect 6419 6762 6559 6810
rect 5839 6758 6559 6762
rect 6611 6758 7196 6810
rect 5562 6752 7196 6758
rect 5562 6750 5981 6752
rect 5562 6698 5595 6750
rect 5647 6746 5981 6750
rect 5647 6698 5787 6746
rect 5562 6694 5787 6698
rect 5839 6700 5981 6746
rect 6033 6750 7196 6752
rect 6033 6700 6173 6750
rect 5839 6698 6173 6700
rect 6225 6698 6367 6750
rect 6419 6746 7196 6750
rect 6419 6698 6559 6746
rect 5839 6694 6559 6698
rect 6611 6694 7196 6746
rect 7970 6779 8114 6802
rect 7970 6727 7984 6779
rect 8036 6727 8048 6779
rect 8100 6727 8114 6779
rect 7970 6704 8114 6727
rect 9952 6720 10044 6734
rect 5562 6688 7196 6694
rect 5562 6686 5981 6688
rect 5562 6634 5595 6686
rect 5647 6682 5981 6686
rect 5647 6634 5787 6682
rect 5562 6630 5787 6634
rect 5839 6636 5981 6682
rect 6033 6686 7196 6688
rect 6033 6636 6173 6686
rect 5839 6634 6173 6636
rect 6225 6634 6367 6686
rect 6419 6684 7196 6686
rect 6419 6682 6624 6684
rect 6419 6634 6559 6682
rect 5839 6630 6559 6634
rect 6611 6630 6624 6682
rect 5562 6626 6624 6630
rect 5592 6614 5650 6626
rect 5784 6610 5842 6626
rect 5978 6616 6036 6626
rect 6170 6614 6228 6626
rect 6364 6614 6422 6626
rect 6556 6610 6614 6626
rect 4626 6457 4902 6498
rect 4626 6085 4642 6457
rect 4886 6085 4902 6457
rect 4626 6044 4902 6085
rect 5688 5962 5746 5976
rect 5688 5948 5691 5962
rect 5654 5934 5691 5948
rect 5332 5910 5691 5934
rect 5743 5948 5746 5962
rect 5882 5966 5940 5986
rect 5882 5948 5885 5966
rect 5743 5914 5885 5948
rect 5937 5948 5940 5966
rect 6074 5964 6132 5984
rect 6074 5948 6077 5964
rect 5937 5914 6077 5948
rect 5743 5912 6077 5914
rect 6129 5948 6132 5964
rect 6266 5950 6324 5970
rect 6266 5948 6269 5950
rect 6129 5912 6269 5948
rect 5743 5910 6269 5912
rect 5332 5902 6269 5910
rect 5332 5898 5885 5902
rect 5332 5846 5691 5898
rect 5743 5850 5885 5898
rect 5937 5900 6269 5902
rect 5937 5850 6077 5900
rect 5743 5848 6077 5850
rect 6129 5898 6269 5900
rect 6321 5948 6324 5950
rect 6458 5950 6516 5970
rect 6458 5948 6461 5950
rect 6321 5898 6461 5948
rect 6513 5948 6516 5950
rect 6513 5898 6540 5948
rect 6129 5886 6540 5898
rect 6129 5848 6269 5886
rect 5743 5846 6269 5848
rect 5332 5838 6269 5846
rect 5332 5832 5885 5838
rect 5332 5780 5473 5832
rect 5525 5786 5885 5832
rect 5937 5836 6269 5838
rect 5937 5786 6077 5836
rect 5525 5784 6077 5786
rect 6129 5834 6269 5836
rect 6321 5834 6461 5886
rect 6513 5834 6540 5886
rect 6129 5822 6540 5834
rect 6129 5784 6269 5822
rect 5525 5780 6269 5784
rect 5332 5774 6269 5780
rect 5332 5768 5885 5774
rect 5332 5716 5473 5768
rect 5525 5722 5885 5768
rect 5937 5772 6269 5774
rect 5937 5722 6077 5772
rect 5525 5720 6077 5722
rect 6129 5770 6269 5772
rect 6321 5770 6461 5822
rect 6513 5770 6540 5822
rect 6129 5758 6540 5770
rect 6129 5720 6269 5758
rect 5525 5716 6269 5720
rect 5332 5710 6269 5716
rect 5332 5704 5885 5710
rect 5332 5652 5473 5704
rect 5525 5658 5885 5704
rect 5937 5708 6269 5710
rect 5937 5658 6077 5708
rect 5525 5656 6077 5658
rect 6129 5706 6269 5708
rect 6321 5706 6461 5758
rect 6513 5706 6540 5758
rect 6129 5694 6540 5706
rect 6129 5656 6269 5694
rect 5525 5652 6269 5656
rect 5332 5646 6269 5652
rect 5332 5638 5885 5646
rect 5332 5632 5691 5638
rect 5654 5586 5691 5632
rect 5743 5594 5885 5638
rect 5937 5644 6269 5646
rect 5937 5594 6077 5644
rect 5743 5592 6077 5594
rect 6129 5642 6269 5644
rect 6321 5642 6461 5694
rect 6513 5642 6540 5694
rect 6129 5630 6540 5642
rect 6129 5592 6269 5630
rect 5743 5586 6269 5592
rect 5654 5582 6269 5586
rect 5654 5574 5885 5582
rect 5654 5522 5691 5574
rect 5743 5530 5885 5574
rect 5937 5580 6269 5582
rect 5937 5530 6077 5580
rect 5743 5528 6077 5530
rect 6129 5578 6269 5580
rect 6321 5578 6461 5630
rect 6513 5578 6540 5630
rect 6129 5566 6540 5578
rect 6129 5528 6269 5566
rect 5743 5522 6269 5528
rect 5654 5514 6269 5522
rect 6321 5514 6461 5566
rect 6513 5514 6540 5566
rect 5688 5500 5746 5514
rect 5882 5510 5940 5514
rect 6074 5508 6132 5514
rect 6266 5494 6324 5514
rect 6458 5494 6516 5514
rect 4144 5124 4316 5126
rect 4142 5115 4326 5124
rect 4142 4979 4162 5115
rect 4298 4979 4326 5115
rect 4142 4974 4326 4979
rect 7074 4986 7194 6684
rect 9952 6664 9970 6720
rect 10026 6664 10044 6720
rect 9952 6650 10044 6664
rect 10344 6542 10482 6558
rect 10344 6486 10345 6542
rect 10401 6540 10425 6542
rect 10407 6488 10419 6540
rect 10401 6486 10425 6488
rect 10481 6486 10482 6542
rect 10344 6470 10482 6486
rect 8288 6377 8342 6392
rect 8288 6362 8289 6377
rect 8276 6325 8289 6362
rect 8341 6362 8342 6377
rect 8480 6377 8534 6392
rect 8480 6362 8481 6377
rect 8341 6333 8481 6362
rect 8533 6362 8534 6377
rect 8684 6362 8760 6364
rect 8533 6344 8770 6362
rect 8533 6333 8696 6344
rect 8341 6325 8478 6333
rect 8276 6313 8478 6325
rect 8276 6276 8289 6313
rect 8288 6261 8289 6276
rect 8341 6277 8478 6313
rect 8534 6292 8696 6333
rect 8748 6292 8770 6344
rect 8534 6277 8770 6292
rect 8341 6276 8481 6277
rect 8341 6261 8342 6276
rect 8476 6266 8481 6276
rect 8288 6246 8342 6261
rect 8480 6261 8481 6266
rect 8533 6276 8770 6277
rect 8533 6266 8536 6276
rect 8684 6272 8760 6276
rect 8533 6261 8534 6266
rect 8480 6246 8534 6261
rect 7794 6228 7872 6244
rect 7794 6226 7811 6228
rect 7794 6174 7801 6226
rect 7794 6172 7811 6174
rect 7867 6172 7872 6228
rect 7794 6156 7872 6172
rect 10594 6150 10642 6998
rect 10866 6788 10996 6800
rect 10864 6764 10996 6788
rect 10864 6712 10873 6764
rect 10925 6757 10937 6764
rect 10989 6712 10996 6764
rect 10864 6701 10898 6712
rect 10954 6701 10996 6712
rect 10864 6676 10996 6701
rect 10864 6670 10988 6676
rect 7512 6122 7578 6144
rect 7512 6070 7519 6122
rect 7571 6120 7578 6122
rect 8178 6142 8244 6144
rect 8572 6142 8638 6144
rect 10594 6142 10678 6150
rect 8178 6122 8654 6142
rect 10100 6136 12748 6142
rect 10072 6126 10610 6136
rect 10072 6122 10091 6126
rect 8178 6120 8185 6122
rect 7571 6070 8185 6120
rect 8237 6120 8579 6122
rect 8237 6070 8383 6120
rect 7512 6068 8383 6070
rect 8435 6070 8579 6120
rect 8631 6070 8654 6122
rect 9884 6120 10091 6122
rect 9874 6118 10091 6120
rect 9868 6074 10091 6118
rect 10143 6084 10610 6126
rect 10662 6126 12748 6136
rect 10662 6120 12668 6126
rect 10662 6084 11126 6120
rect 10143 6074 11126 6084
rect 9868 6072 11126 6074
rect 8435 6068 8654 6070
rect 7512 6042 8654 6068
rect 9378 6057 9444 6072
rect 9378 6054 9385 6057
rect 7512 6040 8244 6042
rect 7578 6020 8178 6040
rect 8376 6038 8442 6042
rect 8572 6040 8638 6042
rect 9378 5998 9381 6054
rect 9437 5998 9444 6057
rect 9378 5990 9444 5998
rect 9868 6062 10610 6072
rect 9868 6010 10091 6062
rect 10143 6020 10610 6062
rect 10662 6068 11126 6072
rect 11178 6112 12668 6120
rect 11178 6068 11644 6112
rect 10662 6060 11644 6068
rect 11696 6060 12156 6112
rect 12208 6074 12668 6112
rect 12720 6074 12748 6126
rect 12208 6062 12748 6074
rect 12208 6060 12668 6062
rect 10662 6056 12668 6060
rect 10662 6020 11126 6056
rect 10143 6010 11126 6020
rect 9868 6008 11126 6010
rect 9868 5998 10610 6008
rect 9380 5988 9438 5990
rect 9868 5946 10091 5998
rect 10143 5956 10610 5998
rect 10662 6004 11126 6008
rect 11178 6048 12668 6056
rect 11178 6004 11644 6048
rect 10662 5996 11644 6004
rect 11696 5996 12156 6048
rect 12208 6010 12668 6048
rect 12720 6010 12748 6062
rect 12208 5998 12748 6010
rect 12208 5996 12668 5998
rect 10662 5992 12668 5996
rect 10662 5956 11126 5992
rect 10143 5946 11126 5956
rect 9868 5944 11126 5946
rect 9114 5930 9166 5942
rect 9868 5934 10610 5944
rect 9868 5930 10091 5934
rect 9114 5926 10091 5930
rect 9166 5882 10091 5926
rect 10143 5892 10610 5934
rect 10662 5940 11126 5944
rect 11178 5984 12668 5992
rect 11178 5940 11644 5984
rect 10662 5932 11644 5940
rect 11696 5932 12156 5984
rect 12208 5946 12668 5984
rect 12720 5946 12748 5998
rect 12208 5934 12748 5946
rect 12208 5932 12668 5934
rect 10662 5928 12668 5932
rect 10662 5892 11126 5928
rect 10143 5882 11126 5892
rect 9166 5880 11126 5882
rect 9868 5878 11126 5880
rect 9868 5876 10226 5878
rect 9884 5874 10226 5876
rect 11110 5876 11126 5878
rect 11178 5920 12668 5928
rect 11178 5878 11644 5920
rect 11178 5876 11194 5878
rect 9114 5858 9166 5874
rect 10072 5872 10162 5874
rect 11110 5862 11194 5876
rect 11628 5868 11644 5878
rect 11696 5878 12156 5920
rect 11696 5868 11712 5878
rect 11628 5854 11712 5868
rect 12140 5868 12156 5878
rect 12208 5882 12668 5920
rect 12720 5882 12748 5934
rect 12208 5878 12748 5882
rect 12208 5868 12224 5878
rect 12652 5868 12736 5878
rect 12140 5854 12224 5868
rect 9024 5722 9202 5736
rect 9024 5666 9045 5722
rect 9101 5720 9125 5722
rect 9107 5668 9119 5720
rect 9101 5666 9125 5668
rect 9181 5666 9202 5722
rect 9024 5652 9202 5666
rect 7904 5385 8122 5408
rect 7904 5363 7923 5385
rect 8103 5363 8122 5385
rect 7904 5227 7905 5363
rect 8121 5227 8122 5363
rect 7904 5205 7923 5227
rect 8103 5205 8122 5227
rect 7904 5182 8122 5205
rect 10332 5134 10408 5188
rect 10846 5134 10950 5152
rect 11370 5134 11474 5138
rect 11874 5134 11978 5148
rect 12392 5136 12496 5152
rect 12290 5134 12600 5136
rect 10270 5127 12604 5134
rect 10270 5122 10872 5127
rect 10246 5113 10872 5122
rect 10246 5091 10352 5113
rect 10404 5091 10872 5113
rect 10246 5035 10350 5091
rect 10406 5075 10872 5091
rect 10924 5123 12418 5127
rect 10924 5113 11900 5123
rect 10924 5075 11396 5113
rect 10406 5063 11396 5075
rect 10406 5035 10872 5063
rect 10246 5011 10352 5035
rect 10404 5011 10872 5035
rect 10924 5061 11396 5063
rect 11448 5071 11900 5113
rect 11952 5075 12418 5123
rect 12470 5075 12604 5127
rect 11952 5071 12604 5075
rect 11448 5063 12604 5071
rect 11448 5061 12418 5063
rect 10924 5059 12418 5061
rect 10924 5049 11900 5059
rect 10924 5011 11396 5049
rect 4144 4968 4316 4974
rect 6034 4868 6098 4888
rect 6034 4858 6038 4868
rect 6034 4806 6037 4858
rect 6094 4812 6098 4868
rect 6089 4806 6098 4812
rect 6034 4792 6098 4806
rect 6146 4866 6216 4878
rect 6146 4860 6153 4866
rect 6146 4808 6149 4860
rect 6209 4810 6216 4866
rect 6201 4808 6216 4810
rect 6146 4798 6216 4808
rect 6146 4796 6204 4798
rect 7074 4760 7218 4986
rect 10246 4955 10350 5011
rect 10406 4999 11396 5011
rect 10406 4955 10872 4999
rect 10246 4933 10352 4955
rect 10404 4947 10872 4955
rect 10924 4997 11396 4999
rect 11448 5007 11900 5049
rect 11952 5011 12418 5059
rect 12470 5011 12604 5063
rect 11952 5007 12604 5011
rect 11448 4999 12604 5007
rect 11448 4997 12418 4999
rect 10924 4995 12418 4997
rect 10924 4985 11900 4995
rect 10924 4947 11396 4985
rect 10404 4933 11396 4947
rect 11448 4943 11900 4985
rect 11952 4947 12418 4995
rect 12470 4947 12604 4999
rect 11952 4943 12604 4947
rect 11448 4933 12604 4943
rect 10246 4930 12604 4933
rect 10270 4920 12604 4930
rect 10340 4914 10416 4920
rect 11370 4908 11474 4920
rect 11874 4918 11978 4920
rect 12290 4878 12600 4920
rect 5922 4738 7218 4760
rect 5922 4686 5929 4738
rect 5981 4686 7218 4738
rect 5922 4678 7218 4686
rect 5922 4672 7210 4678
rect 4230 4543 4304 4562
rect 4230 4487 4241 4543
rect 4297 4487 4304 4543
rect 4230 4464 4304 4487
<< via2 >>
rect 6782 10761 6800 10897
rect 6800 10761 6980 10897
rect 6980 10761 6998 10897
rect 4869 9953 5085 10320
rect 6565 10251 6613 10276
rect 6613 10251 6621 10276
rect 6565 10239 6621 10251
rect 6565 10220 6613 10239
rect 6613 10220 6621 10239
rect 6565 10187 6613 10196
rect 6613 10187 6621 10196
rect 6565 10175 6621 10187
rect 6565 10140 6613 10175
rect 6613 10140 6621 10175
rect 6689 10249 6745 10268
rect 6689 10212 6728 10249
rect 6728 10212 6745 10249
rect 6689 10185 6745 10188
rect 6689 10133 6728 10185
rect 6728 10133 6745 10185
rect 6689 10132 6745 10133
rect 4869 9944 5085 9953
rect 11640 9841 11856 9849
rect 10362 9636 10418 9638
rect 10362 9584 10364 9636
rect 10364 9584 10416 9636
rect 10416 9584 10418 9636
rect 10362 9582 10418 9584
rect 8106 8945 8162 8999
rect 8106 8943 8152 8945
rect 8152 8943 8162 8945
rect 8106 8893 8152 8919
rect 8152 8893 8162 8919
rect 8106 8863 8162 8893
rect 11640 9473 11856 9841
rect 9847 9410 9903 9415
rect 9847 9359 9849 9410
rect 9849 9359 9901 9410
rect 9901 9359 9903 9410
rect 11639 9201 11855 9203
rect 11639 8829 11855 9201
rect 11639 8827 11855 8829
rect 7885 8258 7941 8260
rect 7885 8206 7887 8258
rect 7887 8206 7939 8258
rect 7939 8206 7941 8258
rect 7885 8204 7941 8206
rect 14294 7845 14338 7896
rect 14338 7845 14350 7896
rect 14294 7840 14350 7845
rect 10905 7310 10961 7313
rect 9974 7257 10030 7259
rect 9974 7205 9976 7257
rect 9976 7205 10028 7257
rect 10028 7205 10030 7257
rect 9974 7203 10030 7205
rect 10905 7258 10947 7310
rect 10947 7258 10961 7310
rect 10905 7257 10961 7258
rect 8079 7113 8135 7121
rect 8079 7065 8131 7113
rect 8131 7065 8135 7113
rect 8079 6997 8131 7041
rect 8131 6997 8135 7041
rect 8079 6985 8135 6997
rect 8896 7092 8898 7114
rect 8898 7092 8950 7114
rect 8950 7092 8952 7114
rect 8896 7080 8952 7092
rect 8896 7058 8898 7080
rect 8898 7058 8950 7080
rect 8950 7058 8952 7080
rect 4162 5100 4298 5115
rect 4162 5048 4243 5100
rect 4243 5048 4295 5100
rect 4295 5048 4298 5100
rect 4162 4979 4298 5048
rect 9970 6718 10026 6720
rect 9970 6666 9972 6718
rect 9972 6666 10024 6718
rect 10024 6666 10026 6718
rect 9970 6664 10026 6666
rect 10345 6540 10401 6542
rect 10425 6540 10481 6542
rect 10345 6488 10355 6540
rect 10355 6488 10401 6540
rect 10425 6488 10471 6540
rect 10471 6488 10481 6540
rect 10345 6486 10401 6488
rect 10425 6486 10481 6488
rect 8478 6325 8481 6333
rect 8481 6325 8533 6333
rect 8533 6325 8534 6333
rect 8478 6313 8534 6325
rect 8478 6277 8481 6313
rect 8481 6277 8533 6313
rect 8533 6277 8534 6313
rect 7811 6226 7867 6228
rect 7811 6174 7853 6226
rect 7853 6174 7867 6226
rect 7811 6172 7867 6174
rect 10898 6712 10925 6757
rect 10925 6712 10937 6757
rect 10937 6712 10954 6757
rect 10898 6701 10954 6712
rect 9381 6005 9385 6054
rect 9385 6005 9437 6054
rect 9381 5998 9437 6005
rect 9045 5720 9101 5722
rect 9125 5720 9181 5722
rect 9045 5668 9055 5720
rect 9055 5668 9101 5720
rect 9125 5668 9171 5720
rect 9171 5668 9181 5720
rect 9045 5666 9101 5668
rect 9125 5666 9181 5668
rect 7905 5227 7923 5363
rect 7923 5227 8103 5363
rect 8103 5227 8121 5363
rect 10350 5061 10352 5091
rect 10352 5061 10404 5091
rect 10404 5061 10406 5091
rect 10350 5049 10406 5061
rect 10350 5035 10352 5049
rect 10352 5035 10404 5049
rect 10404 5035 10406 5049
rect 6038 4858 6094 4868
rect 6038 4812 6089 4858
rect 6089 4812 6094 4858
rect 6153 4860 6209 4866
rect 6153 4810 6201 4860
rect 6201 4810 6209 4860
rect 10350 4997 10352 5011
rect 10352 4997 10404 5011
rect 10404 4997 10406 5011
rect 10350 4985 10406 4997
rect 10350 4955 10352 4985
rect 10352 4955 10404 4985
rect 10404 4955 10406 4985
rect 4241 4539 4297 4543
rect 4241 4487 4293 4539
rect 4293 4487 4297 4539
<< metal3 >>
rect 6772 10901 7008 10941
rect 6772 10897 6818 10901
rect 6962 10897 7008 10901
rect 6772 10761 6782 10897
rect 6998 10761 7008 10897
rect 6772 10757 6818 10761
rect 6962 10757 7008 10761
rect 6772 10717 7008 10757
rect 4848 10320 5106 10325
rect 4848 10284 4869 10320
rect 5085 10284 5106 10320
rect 4848 9980 4865 10284
rect 5089 9980 5106 10284
rect 6548 10294 6638 10295
rect 6548 10287 6750 10294
rect 6548 10280 6762 10287
rect 6548 10216 6561 10280
rect 6625 10272 6762 10280
rect 6625 10216 6685 10272
rect 6548 10208 6685 10216
rect 6749 10208 6762 10272
rect 6548 10200 6762 10208
rect 6548 10136 6561 10200
rect 6625 10192 6762 10200
rect 6625 10136 6685 10192
rect 6548 10128 6685 10136
rect 6749 10128 6762 10192
rect 6548 10121 6762 10128
rect 6558 10113 6762 10121
rect 6558 10106 6750 10113
rect 4848 9944 4869 9980
rect 5085 9944 5106 9980
rect 4848 9939 5106 9944
rect 11612 9853 11884 9873
rect 10346 9642 10434 9665
rect 10346 9578 10358 9642
rect 10422 9578 10434 9642
rect 10346 9555 10434 9578
rect 11612 9469 11636 9853
rect 11860 9469 11884 9853
rect 9828 9419 9922 9455
rect 11612 9449 11884 9469
rect 9828 9355 9843 9419
rect 9907 9355 9922 9419
rect 9828 9319 9922 9355
rect 11606 9223 11910 9228
rect 11596 9203 11910 9223
rect 8090 9007 8184 9020
rect 8086 8999 8184 9007
rect 8086 8943 8106 8999
rect 8162 8943 8184 8999
rect 8086 8919 8184 8943
rect 8086 8863 8106 8919
rect 8162 8863 8184 8919
rect 8086 8855 8184 8863
rect 8090 8676 8184 8855
rect 11596 8827 11639 9203
rect 11855 8827 11910 9203
rect 11596 8807 11910 8827
rect 11606 8676 11910 8807
rect 8088 8476 11948 8676
rect 7050 8324 7444 8436
rect 7050 8260 7968 8324
rect 7050 8204 7885 8260
rect 7941 8204 7968 8260
rect 7050 8128 7968 8204
rect 4134 5115 4326 5121
rect 4134 5079 4162 5115
rect 4298 5079 4326 5115
rect 4134 5015 4158 5079
rect 4302 5015 4326 5079
rect 4134 4979 4162 5015
rect 4298 4979 4326 5015
rect 4134 4973 4326 4979
rect 6024 4882 6108 4883
rect 7050 4882 7444 8128
rect 14282 7903 14380 7920
rect 14282 7896 14299 7903
rect 14282 7840 14294 7896
rect 14282 7839 14299 7840
rect 14363 7839 14380 7903
rect 14282 7822 14380 7839
rect 14282 7817 14362 7822
rect 10866 7317 11000 7337
rect 9950 7263 10054 7281
rect 8894 7168 9006 7206
rect 9950 7199 9970 7263
rect 10034 7199 10054 7263
rect 10866 7253 10901 7317
rect 10965 7253 11000 7317
rect 10866 7233 11000 7253
rect 9950 7181 10054 7199
rect 8884 7148 9006 7168
rect 8052 7125 8162 7143
rect 8052 7061 8075 7125
rect 8139 7061 8162 7125
rect 8052 7045 8162 7061
rect 8052 6981 8075 7045
rect 8139 6981 8162 7045
rect 8052 6963 8162 6981
rect 8882 7140 9006 7148
rect 8882 7114 8998 7140
rect 8882 7058 8896 7114
rect 8952 7066 8998 7114
rect 8952 7058 9004 7066
rect 8882 6976 9004 7058
rect 7792 6232 7914 6846
rect 7792 6168 7807 6232
rect 7871 6168 7914 6232
rect 7792 6144 7914 6168
rect 8464 6333 8556 6386
rect 8464 6277 8478 6333
rect 8534 6277 8556 6333
rect 7894 5396 8132 5403
rect 7854 5363 8136 5396
rect 7854 5227 7905 5363
rect 8121 5354 8136 5363
rect 8464 5354 8556 6277
rect 8882 5732 8970 6976
rect 10856 6784 10988 6798
rect 10856 6783 11008 6784
rect 9938 6736 10070 6760
rect 10854 6757 11008 6783
rect 10854 6736 10898 6757
rect 9938 6720 10898 6736
rect 9938 6664 9970 6720
rect 10026 6701 10898 6720
rect 10954 6701 11008 6757
rect 10026 6676 11008 6701
rect 10026 6672 11004 6676
rect 10026 6664 10988 6672
rect 9938 6660 10988 6664
rect 9942 6655 10988 6660
rect 9944 6654 10988 6655
rect 9958 6642 10984 6654
rect 10334 6546 10492 6553
rect 10334 6542 10381 6546
rect 10445 6542 10492 6546
rect 10334 6486 10345 6542
rect 10481 6486 10492 6542
rect 10334 6482 10381 6486
rect 10445 6482 10492 6486
rect 10334 6475 10492 6482
rect 9376 6059 9468 6062
rect 9370 6054 9468 6059
rect 9370 5998 9381 6054
rect 9437 5998 9468 6054
rect 9370 5993 9468 5998
rect 9376 5946 9468 5993
rect 8882 5731 9102 5732
rect 8882 5722 9212 5731
rect 8882 5666 9045 5722
rect 9101 5666 9125 5722
rect 9181 5666 9212 5722
rect 8882 5657 9212 5666
rect 8882 5598 9162 5657
rect 8882 5354 8970 5598
rect 9400 5354 9468 5946
rect 8121 5334 9178 5354
rect 9340 5334 9486 5354
rect 8121 5227 9486 5334
rect 7854 5204 9486 5227
rect 7854 4882 8136 5204
rect 8882 5178 8970 5204
rect 9102 5200 9422 5204
rect 10332 5127 10408 5188
rect 10330 5095 10426 5127
rect 10330 5031 10346 5095
rect 10410 5031 10426 5095
rect 10330 5015 10426 5031
rect 10330 4951 10346 5015
rect 10410 4951 10426 5015
rect 10330 4919 10426 4951
rect 6024 4868 8162 4882
rect 6024 4812 6038 4868
rect 6094 4866 8162 4868
rect 6094 4812 6153 4866
rect 6024 4810 6153 4812
rect 6209 4810 8162 4866
rect 6024 4802 8162 4810
rect 6024 4797 6108 4802
rect 4198 4543 4314 4566
rect 4198 4487 4241 4543
rect 4297 4487 4314 4543
rect 4198 4444 4314 4487
rect 7050 4444 7444 4802
rect 7854 4444 8136 4802
rect 4178 4242 8192 4444
rect 4590 4240 5020 4242
rect 7050 4238 7444 4242
rect 7854 4220 8136 4242
<< via3 >>
rect 6818 10897 6962 10901
rect 6818 10761 6962 10897
rect 6818 10757 6962 10761
rect 4865 9980 4869 10284
rect 4869 9980 5085 10284
rect 5085 9980 5089 10284
rect 6561 10276 6625 10280
rect 6561 10220 6565 10276
rect 6565 10220 6621 10276
rect 6621 10220 6625 10276
rect 6561 10216 6625 10220
rect 6685 10268 6749 10272
rect 6685 10212 6689 10268
rect 6689 10212 6745 10268
rect 6745 10212 6749 10268
rect 6685 10208 6749 10212
rect 6561 10196 6625 10200
rect 6561 10140 6565 10196
rect 6565 10140 6621 10196
rect 6621 10140 6625 10196
rect 6561 10136 6625 10140
rect 6685 10188 6749 10192
rect 6685 10132 6689 10188
rect 6689 10132 6745 10188
rect 6745 10132 6749 10188
rect 6685 10128 6749 10132
rect 10358 9638 10422 9642
rect 10358 9582 10362 9638
rect 10362 9582 10418 9638
rect 10418 9582 10422 9638
rect 10358 9578 10422 9582
rect 11636 9849 11860 9853
rect 11636 9473 11640 9849
rect 11640 9473 11856 9849
rect 11856 9473 11860 9849
rect 11636 9469 11860 9473
rect 9843 9415 9907 9419
rect 9843 9359 9847 9415
rect 9847 9359 9903 9415
rect 9903 9359 9907 9415
rect 9843 9355 9907 9359
rect 4158 5015 4162 5079
rect 4162 5015 4222 5079
rect 4238 5015 4298 5079
rect 4298 5015 4302 5079
rect 14299 7896 14363 7903
rect 14299 7840 14350 7896
rect 14350 7840 14363 7896
rect 14299 7839 14363 7840
rect 9970 7259 10034 7263
rect 9970 7203 9974 7259
rect 9974 7203 10030 7259
rect 10030 7203 10034 7259
rect 9970 7199 10034 7203
rect 10901 7313 10965 7317
rect 10901 7257 10905 7313
rect 10905 7257 10961 7313
rect 10961 7257 10965 7313
rect 10901 7253 10965 7257
rect 8075 7121 8139 7125
rect 8075 7065 8079 7121
rect 8079 7065 8135 7121
rect 8135 7065 8139 7121
rect 8075 7061 8139 7065
rect 8075 7041 8139 7045
rect 8075 6985 8079 7041
rect 8079 6985 8135 7041
rect 8135 6985 8139 7041
rect 8075 6981 8139 6985
rect 7807 6228 7871 6232
rect 7807 6172 7811 6228
rect 7811 6172 7867 6228
rect 7867 6172 7871 6228
rect 7807 6168 7871 6172
rect 10381 6542 10445 6546
rect 10381 6486 10401 6542
rect 10401 6486 10425 6542
rect 10425 6486 10445 6542
rect 10381 6482 10445 6486
rect 10346 5091 10410 5095
rect 10346 5035 10350 5091
rect 10350 5035 10406 5091
rect 10406 5035 10410 5091
rect 10346 5031 10410 5035
rect 10346 5011 10410 5015
rect 10346 4955 10350 5011
rect 10350 4955 10406 5011
rect 10406 4955 10410 5011
rect 10346 4951 10410 4955
<< metal4 >>
rect 4818 10950 5116 10954
rect 4748 10948 6976 10950
rect 4132 10937 6976 10948
rect 4132 10901 6999 10937
rect 4132 10757 6818 10901
rect 6962 10892 6999 10901
rect 7084 10892 7316 10902
rect 9552 10892 9912 10900
rect 6962 10802 9912 10892
rect 6962 10757 9916 10802
rect 4132 10742 9916 10757
rect 4132 10740 9654 10742
rect 4132 10738 7780 10740
rect 7908 10738 9654 10740
rect 4132 10734 6999 10738
rect 4132 10720 5116 10734
rect 6781 10721 6999 10734
rect 4142 5117 4296 10720
rect 4818 10284 5116 10720
rect 7084 10294 7316 10738
rect 9846 10294 9916 10742
rect 10876 10294 10994 10316
rect 11812 10294 12210 10296
rect 14288 10294 14386 10308
rect 4818 9980 4865 10284
rect 5089 9980 5116 10284
rect 6554 10280 7328 10294
rect 6554 10216 6561 10280
rect 6625 10272 7328 10280
rect 6625 10216 6685 10272
rect 6554 10208 6685 10216
rect 6749 10208 7328 10272
rect 6554 10200 7328 10208
rect 6554 10136 6561 10200
rect 6625 10192 7328 10200
rect 6625 10136 6685 10192
rect 6554 10128 6685 10136
rect 6749 10128 7328 10192
rect 9766 10176 14386 10294
rect 6554 10124 7328 10128
rect 6556 10122 6792 10124
rect 6556 10117 6753 10122
rect 6556 10114 6752 10117
rect 4818 9910 5116 9980
rect 7084 6848 7316 10124
rect 9854 9451 9932 10176
rect 10336 10128 10480 10176
rect 9837 9419 9932 9451
rect 9837 9355 9843 9419
rect 9907 9355 9932 9419
rect 9837 9323 9932 9355
rect 9854 7404 9932 9323
rect 9850 7282 9932 7404
rect 10340 9642 10478 10128
rect 10340 9578 10358 9642
rect 10422 9578 10478 9642
rect 9850 7280 10040 7282
rect 9850 7263 10052 7280
rect 9850 7199 9970 7263
rect 10034 7199 10052 7263
rect 9850 7196 10052 7199
rect 9926 7188 10052 7196
rect 9959 7185 10045 7188
rect 8056 7139 8116 7156
rect 8056 7125 8153 7139
rect 8056 7061 8075 7125
rect 8139 7061 8153 7125
rect 8056 7045 8153 7061
rect 8056 6981 8075 7045
rect 8139 6981 8153 7045
rect 8056 6967 8153 6981
rect 8056 6848 8116 6967
rect 7084 6696 8202 6848
rect 10340 6834 10478 9578
rect 10876 7333 10994 10176
rect 11606 10170 12210 10176
rect 11606 9853 11882 10170
rect 11606 9469 11636 9853
rect 11860 9469 11882 9853
rect 11606 9458 11882 9469
rect 11621 9453 11875 9458
rect 14288 7903 14386 10176
rect 14288 7839 14299 7903
rect 14363 7839 14386 7903
rect 14288 7804 14386 7839
rect 10875 7317 10994 7333
rect 10875 7253 10901 7317
rect 10965 7253 10994 7317
rect 10875 7248 10994 7253
rect 10875 7237 10991 7248
rect 7084 6690 7316 6696
rect 7730 6682 7914 6696
rect 7792 6232 7914 6682
rect 10340 6656 10482 6834
rect 7792 6168 7807 6232
rect 7871 6168 7914 6232
rect 7792 6144 7914 6168
rect 10342 6549 10482 6656
rect 10342 6546 10483 6549
rect 10342 6482 10381 6546
rect 10445 6482 10483 6546
rect 10342 6479 10483 6482
rect 10342 5188 10482 6479
rect 10332 5122 10482 5188
rect 4142 5079 4317 5117
rect 4142 5015 4158 5079
rect 4222 5015 4238 5079
rect 4302 5015 4317 5079
rect 4142 5002 4317 5015
rect 4143 4977 4317 5002
rect 10339 5095 10482 5122
rect 10339 5031 10346 5095
rect 10410 5031 10482 5095
rect 10339 5015 10482 5031
rect 10339 4951 10346 5015
rect 10410 4951 10482 5015
rect 10339 4926 10482 4951
rect 10339 4924 10478 4926
rect 10339 4923 10417 4924
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1724995455
transform 1 0 6017 0 1 4772
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_9B2JY7  sky130_fd_pr__nfet_01v8_9B2JY7_0
timestamp 1724995455
transform 0 -1 11364 1 0 11485
box -349 -1100 349 1100
use sky130_fd_pr__nfet_01v8_U2JGXT  sky130_fd_pr__nfet_01v8_U2JGXT_0
timestamp 1724995455
transform 0 1 8396 -1 0 8206
box -216 -500 216 500
use sky130_fd_pr__res_xhigh_po_1p41_VHK7CU  sky130_fd_pr__res_xhigh_po_1p41_VHK7CU_0
timestamp 1724995455
transform 1 0 11752 0 1 9335
box -297 -694 297 694
use sky130_fd_pr__res_xhigh_po_1p41_VHK7CU  sky130_fd_pr__res_xhigh_po_1p41_VHK7CU_1
timestamp 1724995455
transform 1 0 4959 0 1 9804
box -297 -694 297 694
use sky130_fd_pr__res_xhigh_po_1p41_VHK7CU  sky130_fd_pr__res_xhigh_po_1p41_VHK7CU_2
timestamp 1724995455
transform 1 0 4759 0 1 6622
box -297 -694 297 694
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1724995455
transform 1 0 4070 0 1 4524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1724995455
transform 1 0 10226 0 1 6688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1724995455
transform 1 0 10800 0 1 6696
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1724995455
transform 1 0 4228 0 1 4520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x5
timestamp 1724995455
transform 1 0 10892 0 1 6696
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1724995455
transform 1 0 9958 0 1 6688
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_SKB8VM  XM4
timestamp 1724995455
transform 1 0 6100 0 1 7975
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_SKB8VM  XM5
timestamp 1724995455
transform -1 0 6076 0 -1 9087
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_SKB8VM  XM6
timestamp 1724995455
transform -1 0 6056 0 -1 10179
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_VC5S4W  XM7
timestamp 1724995455
transform -1 0 6103 0 -1 6283
box -647 -1019 647 1019
use sky130_fd_pr__nfet_01v8_69TQ3K  XM8
timestamp 1724995455
transform 1 0 9268 0 1 5966
box -286 -300 286 300
use sky130_fd_pr__pfet_01v8_UGNVTG  XM9
timestamp 1724995455
transform -1 0 7809 0 -1 9641
box -359 -1119 359 1119
use sky130_fd_pr__pfet_01v8_XGS3BL  XM10
timestamp 1724995455
transform 1 0 10019 0 1 9509
box -407 -419 407 419
use sky130_fd_pr__nfet_01v8_MSLS59  XM11
timestamp 1724995455
transform 1 0 8407 0 1 6088
box -349 -500 349 500
use sky130_fd_pr__pfet_01v8_3HMWVM  XM12
timestamp 1724995455
transform 1 0 7684 0 1 6149
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_PDPE9S  XM13
timestamp 1724995455
transform 1 0 11409 0 1 5529
box -1457 -1019 1457 1019
use sky130_fd_pr__nfet_01v8_SC2JGL  XM14
timestamp 1724995455
transform 1 0 8681 0 1 7192
box -397 -400 397 400
use sky130_fd_pr__pfet_01v8_XGSNAL  XM15
timestamp 1724995455
transform 1 0 8039 0 1 7241
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_KRS3CJ  XM16
timestamp 1724995455
transform 1 0 11784 0 1 7869
box -2696 -319 2696 319
<< labels >>
flabel metal2 s 6786 10732 6986 10932 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 s 7576 7088 7776 7288 0 FreeSans 320 0 0 0 Va
port 2 nsew
flabel metal1 s 4362 7526 4562 7726 0 FreeSans 320 0 0 0 PAD
port 3 nsew
flabel metal1 s 9240 7180 9436 7380 0 FreeSans 320 0 0 0 Vb
port 4 nsew
flabel metal2 s 7904 5192 8104 5392 0 FreeSans 320 0 0 0 VSS
port 5 nsew
flabel metal1 s 11630 7092 11828 7286 0 FreeSans 320 0 0 0 Vout
port 6 nsew
<< end >>
