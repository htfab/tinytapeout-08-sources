magic
tech sky130A
magscale 1 2
timestamp 1724348452
<< viali >>
rect 1160 1640 1398 1692
rect 1096 -1378 1434 -1330
<< metal1 >>
rect 358 1966 1404 2138
rect 358 1882 376 1966
rect 576 1882 1404 1966
rect 376 1760 576 1766
rect 1148 1704 1404 1882
rect 1138 1692 1422 1704
rect 658 1662 858 1666
rect -136 1600 942 1662
rect 1138 1640 1160 1692
rect 1398 1640 1422 1692
rect 1138 1630 1422 1640
rect -136 1590 958 1600
rect -136 1532 1380 1590
rect -136 1526 958 1532
rect -136 1462 942 1526
rect -136 528 64 1462
rect 370 908 376 1108
rect 576 908 1154 1108
rect 1405 837 2510 1171
rect -136 464 942 528
rect -136 394 1378 464
rect -136 328 942 394
rect 2176 351 2510 837
rect -136 206 64 328
rect -682 6 64 206
rect -136 -44 64 6
rect 2176 17 2729 351
rect -136 -116 956 -44
rect -136 -164 1382 -116
rect -136 -244 956 -164
rect -136 -1156 64 -244
rect 2176 -521 2510 17
rect 386 -796 392 -596
rect 592 -796 1154 -596
rect 1389 -855 2510 -521
rect -136 -1228 972 -1156
rect -136 -1280 1376 -1228
rect -136 -1292 976 -1280
rect -136 -1356 972 -1292
rect 1082 -1330 1458 -1316
rect 1082 -1378 1096 -1330
rect 1434 -1378 1458 -1330
rect 392 -1424 592 -1418
rect 1082 -1526 1458 -1378
rect 392 -1656 592 -1624
rect 1198 -1656 1346 -1526
rect 392 -1804 1346 -1656
rect 392 -1806 592 -1804
<< via1 >>
rect 376 1766 576 1966
rect 376 908 576 1108
rect 392 -796 592 -596
rect 392 -1624 592 -1424
<< metal2 >>
rect 370 1766 376 1966
rect 576 1766 582 1966
rect 376 1108 576 1766
rect 376 902 576 908
rect 392 -596 592 -590
rect 392 -1424 592 -796
rect 386 -1624 392 -1424
rect 592 -1624 598 -1424
use sky130_fd_pr__nfet_01v8_MMMA4V  XM1
timestamp 1724342599
transform 1 0 1266 0 1 -700
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM2
timestamp 1724342599
transform 1 0 1272 0 1 997
box -296 -719 296 719
<< labels >>
flabel metal1 -682 6 -482 206 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 376 1920 576 2120 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 392 -1806 592 -1606 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 2274 86 2474 286 0 FreeSans 256 0 0 0 OUT
port 3 nsew
<< end >>
