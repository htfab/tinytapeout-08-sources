** sch_path: tb.sch
**.subckt tb
V1 VGND 0 0
V2 VPWR 0 3.3
x1 0 0 0 VOUT 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 VGND VPWR
+ tt_um_htfab_pi_snake
**** begin user architecture code
.lib ../../pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.include tt_um_htfab_pi_snake.spice

.control
save all
tran 10n 6u
write snake.raw
.endc

**** end user architecture code
**.ends
.end
