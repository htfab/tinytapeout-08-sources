magic
tech sky130A
magscale 1 2
timestamp 1724342599
<< nwell >>
rect -696 -519 696 519
<< pmos >>
rect -500 -300 500 300
<< pdiff >>
rect -558 288 -500 300
rect -558 -288 -546 288
rect -512 -288 -500 288
rect -558 -300 -500 -288
rect 500 288 558 300
rect 500 -288 512 288
rect 546 -288 558 288
rect 500 -300 558 -288
<< pdiffc >>
rect -546 -288 -512 288
rect 512 -288 546 288
<< nsubdiff >>
rect -660 449 -564 483
rect 564 449 660 483
rect -660 387 -626 449
rect 626 387 660 449
rect -660 -449 -626 -387
rect 626 -449 660 -387
rect -660 -483 -564 -449
rect 564 -483 660 -449
<< nsubdiffcont >>
rect -564 449 564 483
rect -660 -387 -626 387
rect 626 -387 660 387
rect -564 -483 564 -449
<< poly >>
rect -500 381 500 397
rect -500 347 -484 381
rect 484 347 500 381
rect -500 300 500 347
rect -500 -347 500 -300
rect -500 -381 -484 -347
rect 484 -381 500 -347
rect -500 -397 500 -381
<< polycont >>
rect -484 347 484 381
rect -484 -381 484 -347
<< locali >>
rect -660 449 -564 483
rect 564 449 660 483
rect -660 387 -626 449
rect 626 387 660 449
rect -500 347 -484 381
rect 484 347 500 381
rect -546 288 -512 304
rect -546 -304 -512 -288
rect 512 288 546 304
rect 512 -304 546 -288
rect -500 -381 -484 -347
rect 484 -381 500 -347
rect -660 -449 -626 -387
rect 626 -449 660 -387
rect -660 -483 -564 -449
rect 564 -483 660 -449
<< viali >>
rect -484 347 484 381
rect -546 -288 -512 288
rect 512 -288 546 288
rect -484 -381 484 -347
<< metal1 >>
rect -496 381 496 387
rect -496 347 -484 381
rect 484 347 496 381
rect -496 341 496 347
rect -552 288 -506 300
rect -552 -288 -546 288
rect -512 -288 -506 288
rect -552 -300 -506 -288
rect 506 288 552 300
rect 506 -288 512 288
rect 546 -288 552 288
rect 506 -300 552 -288
rect -496 -347 496 -341
rect -496 -381 -484 -347
rect 484 -381 496 -347
rect -496 -387 496 -381
<< properties >>
string FIXED_BBOX -643 -466 643 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
