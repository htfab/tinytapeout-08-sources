magic
tech sky130A
magscale 1 2
timestamp 1725528192
<< pwell >>
rect -367 -685 367 685
<< psubdiff >>
rect -331 615 331 649
rect -331 553 -297 615
rect 297 553 331 615
rect -331 -615 -297 -553
rect 297 -615 331 -553
rect -331 -649 331 -615
<< psubdiffcont >>
rect -331 -553 -297 553
rect 297 -553 331 553
<< xpolycontact >>
rect -201 87 -131 519
rect -201 -519 -131 -87
rect -35 87 35 519
rect -35 -519 35 -87
rect 131 87 201 519
rect 131 -519 201 -87
<< xpolyres >>
rect -201 -87 -131 87
rect -35 -87 35 87
rect 131 -87 201 87
<< locali >>
rect -331 615 331 649
rect -331 553 -297 615
rect 297 553 331 615
rect -331 -615 -297 -553
rect 297 -615 331 -553
rect -331 -649 331 -615
<< viali >>
rect -185 104 -147 501
rect -19 104 19 501
rect 147 104 185 501
rect -185 -501 -147 -104
rect -19 -501 19 -104
rect 147 -501 185 -104
<< metal1 >>
rect -191 501 -141 513
rect -191 104 -185 501
rect -147 104 -141 501
rect -191 92 -141 104
rect -25 501 25 513
rect -25 104 -19 501
rect 19 104 25 501
rect -25 92 25 104
rect 141 501 191 513
rect 141 104 147 501
rect 185 104 191 501
rect 141 92 191 104
rect -191 -104 -141 -92
rect -191 -501 -185 -104
rect -147 -501 -141 -104
rect -191 -513 -141 -501
rect -25 -104 25 -92
rect -25 -501 -19 -104
rect 19 -501 25 -104
rect -25 -513 25 -501
rect 141 -104 191 -92
rect 141 -501 147 -104
rect 185 -501 191 -104
rect 141 -513 191 -501
<< properties >>
string FIXED_BBOX -314 -632 314 632
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.03 m 1 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 6.961k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
