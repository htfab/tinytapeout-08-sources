magic
tech sky130A
magscale 1 2
timestamp 1724943425
<< nmoslvt >>
rect -366 -169 -266 231
rect -208 -169 -108 231
rect -50 -169 50 231
rect 108 -169 208 231
rect 266 -169 366 231
<< ndiff >>
rect -424 219 -366 231
rect -424 -157 -412 219
rect -378 -157 -366 219
rect -424 -169 -366 -157
rect -266 219 -208 231
rect -266 -157 -254 219
rect -220 -157 -208 219
rect -266 -169 -208 -157
rect -108 219 -50 231
rect -108 -157 -96 219
rect -62 -157 -50 219
rect -108 -169 -50 -157
rect 50 219 108 231
rect 50 -157 62 219
rect 96 -157 108 219
rect 50 -169 108 -157
rect 208 219 266 231
rect 208 -157 220 219
rect 254 -157 266 219
rect 208 -169 266 -157
rect 366 219 424 231
rect 366 -157 378 219
rect 412 -157 424 219
rect 366 -169 424 -157
<< ndiffc >>
rect -412 -157 -378 219
rect -254 -157 -220 219
rect -96 -157 -62 219
rect 62 -157 96 219
rect 220 -157 254 219
rect 378 -157 412 219
<< poly >>
rect -366 231 -266 257
rect -208 231 -108 257
rect -50 231 50 257
rect 108 231 208 257
rect 266 231 366 257
rect -366 -207 -266 -169
rect -366 -241 -350 -207
rect -282 -241 -266 -207
rect -366 -257 -266 -241
rect -208 -207 -108 -169
rect -208 -241 -192 -207
rect -124 -241 -108 -207
rect -208 -257 -108 -241
rect -50 -207 50 -169
rect -50 -241 -34 -207
rect 34 -241 50 -207
rect -50 -257 50 -241
rect 108 -207 208 -169
rect 108 -241 124 -207
rect 192 -241 208 -207
rect 108 -257 208 -241
rect 266 -207 366 -169
rect 266 -241 282 -207
rect 350 -241 366 -207
rect 266 -257 366 -241
<< polycont >>
rect -350 -241 -282 -207
rect -192 -241 -124 -207
rect -34 -241 34 -207
rect 124 -241 192 -207
rect 282 -241 350 -207
<< locali >>
rect -412 219 -378 235
rect -412 -173 -378 -157
rect -254 219 -220 235
rect -254 -173 -220 -157
rect -96 219 -62 235
rect -96 -173 -62 -157
rect 62 219 96 235
rect 62 -173 96 -157
rect 220 219 254 235
rect 220 -173 254 -157
rect 378 219 412 235
rect 378 -173 412 -157
rect -366 -241 -350 -207
rect -282 -241 -266 -207
rect -208 -241 -192 -207
rect -124 -241 -108 -207
rect -50 -241 -34 -207
rect 34 -241 50 -207
rect 108 -241 124 -207
rect 192 -241 208 -207
rect 266 -241 282 -207
rect 350 -241 366 -207
<< viali >>
rect -412 89 -378 202
rect -254 -140 -220 -27
rect -96 89 -62 202
rect 62 -140 96 -27
rect 220 89 254 202
rect 378 -140 412 -27
rect -350 -241 -282 -207
rect -192 -241 -124 -207
rect -34 -241 34 -207
rect 124 -241 192 -207
rect 282 -241 350 -207
<< metal1 >>
rect -418 202 -372 214
rect -418 89 -412 202
rect -378 89 -372 202
rect -418 77 -372 89
rect -102 202 -56 214
rect -102 89 -96 202
rect -62 89 -56 202
rect -102 77 -56 89
rect 214 202 260 214
rect 214 89 220 202
rect 254 89 260 202
rect 214 77 260 89
rect -260 -27 -214 -15
rect -260 -140 -254 -27
rect -220 -140 -214 -27
rect -260 -152 -214 -140
rect 56 -27 102 -15
rect 56 -140 62 -27
rect 96 -140 102 -27
rect 56 -152 102 -140
rect 372 -27 418 -15
rect 372 -140 378 -27
rect 412 -140 418 -27
rect 372 -152 418 -140
rect -362 -207 -270 -201
rect -362 -241 -350 -207
rect -282 -241 -270 -207
rect -362 -247 -270 -241
rect -204 -207 -112 -201
rect -204 -241 -192 -207
rect -124 -241 -112 -207
rect -204 -247 -112 -241
rect -46 -207 46 -201
rect -46 -241 -34 -207
rect 34 -241 46 -207
rect -46 -247 46 -241
rect 112 -207 204 -201
rect 112 -241 124 -207
rect 192 -241 204 -207
rect 112 -247 204 -241
rect 270 -207 362 -201
rect 270 -241 282 -207
rect 350 -241 362 -207
rect 270 -247 362 -241
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
