magic
tech sky130A
magscale 1 2
timestamp 1724420584
<< metal1 >>
rect -23327 10441 -23321 10996
rect -22766 10441 -22760 10996
rect -23321 7538 -22766 10441
rect -5832 10352 -4176 11658
rect -5832 10081 8374 10352
rect -22185 9367 8374 10081
rect -5706 9241 8374 9367
rect 7330 9162 8374 9241
rect 7330 9130 7632 9162
rect 7394 9026 7548 9130
rect 6076 8791 6634 8850
rect -23321 6983 -21753 7538
rect -18401 7184 -17894 7384
rect -14369 7164 -13776 7364
rect -10275 7142 -9694 7342
rect -6204 7122 -5660 7322
rect -2171 7102 -1598 7302
rect 1901 7080 2464 7280
rect 6076 7266 6634 8233
rect 11112 7654 12008 7754
rect 11112 7342 12018 7654
rect 5944 7066 6634 7266
rect 9514 7142 12018 7342
rect 6076 6822 6634 7066
rect 11112 6758 12018 7142
rect 11112 6626 12008 6758
rect -22238 4466 7800 5326
rect -5410 3228 -4028 4466
<< via1 >>
rect -23321 10441 -22766 10996
rect 6076 8233 6634 8791
<< metal2 >>
rect -23321 10996 -22766 11002
rect -7481 10996 6634 10997
rect -22766 10441 6634 10996
rect -23321 10435 -22766 10441
rect -7481 10439 6634 10441
rect 6076 8791 6634 10439
rect 6070 8233 6076 8791
rect 6634 8233 6640 8791
use not1  x1
timestamp 1724347750
transform 1 0 -21625 0 1 7036
box -643 -1920 3424 2729
use not1  x2
timestamp 1724347750
transform 1 0 -17593 0 1 7016
box -643 -1920 3424 2729
use not1  x3
timestamp 1724347750
transform 1 0 -13499 0 1 6994
box -643 -1920 3424 2729
use not1  x4
timestamp 1724347750
transform 1 0 -9427 0 1 6974
box -643 -1920 3424 2729
use not1  x5
timestamp 1724347750
transform 1 0 -5395 0 1 6954
box -643 -1920 3424 2729
use not1  x6
timestamp 1724347750
transform 1 0 -1323 0 1 6932
box -643 -1920 3424 2729
use not1  x7
timestamp 1724347750
transform 1 0 2733 0 1 6918
box -643 -1920 3424 2729
use notbig  x8
timestamp 1724348452
transform 1 0 6972 0 1 7060
box -682 -1806 2729 2138
<< labels >>
flabel metal1 -5056 10318 -4856 10518 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 11380 7142 11580 7342 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 -4930 3700 -4730 3900 0 FreeSans 256 0 0 0 VSS
port 2 nsew
<< end >>
