magic
tech sky130A
magscale 1 2
timestamp 1725402679
<< nwell >>
rect -1803 -598 1803 564
<< pmoslvt >>
rect -1709 -536 -1609 464
rect -1551 -536 -1451 464
rect -1393 -536 -1293 464
rect -1235 -536 -1135 464
rect -1077 -536 -977 464
rect -919 -536 -819 464
rect -761 -536 -661 464
rect -603 -536 -503 464
rect -445 -536 -345 464
rect -287 -536 -187 464
rect -129 -536 -29 464
rect 29 -536 129 464
rect 187 -536 287 464
rect 345 -536 445 464
rect 503 -536 603 464
rect 661 -536 761 464
rect 819 -536 919 464
rect 977 -536 1077 464
rect 1135 -536 1235 464
rect 1293 -536 1393 464
rect 1451 -536 1551 464
rect 1609 -536 1709 464
<< pdiff >>
rect -1767 452 -1709 464
rect -1767 -524 -1755 452
rect -1721 -524 -1709 452
rect -1767 -536 -1709 -524
rect -1609 452 -1551 464
rect -1609 -524 -1597 452
rect -1563 -524 -1551 452
rect -1609 -536 -1551 -524
rect -1451 452 -1393 464
rect -1451 -524 -1439 452
rect -1405 -524 -1393 452
rect -1451 -536 -1393 -524
rect -1293 452 -1235 464
rect -1293 -524 -1281 452
rect -1247 -524 -1235 452
rect -1293 -536 -1235 -524
rect -1135 452 -1077 464
rect -1135 -524 -1123 452
rect -1089 -524 -1077 452
rect -1135 -536 -1077 -524
rect -977 452 -919 464
rect -977 -524 -965 452
rect -931 -524 -919 452
rect -977 -536 -919 -524
rect -819 452 -761 464
rect -819 -524 -807 452
rect -773 -524 -761 452
rect -819 -536 -761 -524
rect -661 452 -603 464
rect -661 -524 -649 452
rect -615 -524 -603 452
rect -661 -536 -603 -524
rect -503 452 -445 464
rect -503 -524 -491 452
rect -457 -524 -445 452
rect -503 -536 -445 -524
rect -345 452 -287 464
rect -345 -524 -333 452
rect -299 -524 -287 452
rect -345 -536 -287 -524
rect -187 452 -129 464
rect -187 -524 -175 452
rect -141 -524 -129 452
rect -187 -536 -129 -524
rect -29 452 29 464
rect -29 -524 -17 452
rect 17 -524 29 452
rect -29 -536 29 -524
rect 129 452 187 464
rect 129 -524 141 452
rect 175 -524 187 452
rect 129 -536 187 -524
rect 287 452 345 464
rect 287 -524 299 452
rect 333 -524 345 452
rect 287 -536 345 -524
rect 445 452 503 464
rect 445 -524 457 452
rect 491 -524 503 452
rect 445 -536 503 -524
rect 603 452 661 464
rect 603 -524 615 452
rect 649 -524 661 452
rect 603 -536 661 -524
rect 761 452 819 464
rect 761 -524 773 452
rect 807 -524 819 452
rect 761 -536 819 -524
rect 919 452 977 464
rect 919 -524 931 452
rect 965 -524 977 452
rect 919 -536 977 -524
rect 1077 452 1135 464
rect 1077 -524 1089 452
rect 1123 -524 1135 452
rect 1077 -536 1135 -524
rect 1235 452 1293 464
rect 1235 -524 1247 452
rect 1281 -524 1293 452
rect 1235 -536 1293 -524
rect 1393 452 1451 464
rect 1393 -524 1405 452
rect 1439 -524 1451 452
rect 1393 -536 1451 -524
rect 1551 452 1609 464
rect 1551 -524 1563 452
rect 1597 -524 1609 452
rect 1551 -536 1609 -524
rect 1709 452 1767 464
rect 1709 -524 1721 452
rect 1755 -524 1767 452
rect 1709 -536 1767 -524
<< pdiffc >>
rect -1755 -524 -1721 452
rect -1597 -524 -1563 452
rect -1439 -524 -1405 452
rect -1281 -524 -1247 452
rect -1123 -524 -1089 452
rect -965 -524 -931 452
rect -807 -524 -773 452
rect -649 -524 -615 452
rect -491 -524 -457 452
rect -333 -524 -299 452
rect -175 -524 -141 452
rect -17 -524 17 452
rect 141 -524 175 452
rect 299 -524 333 452
rect 457 -524 491 452
rect 615 -524 649 452
rect 773 -524 807 452
rect 931 -524 965 452
rect 1089 -524 1123 452
rect 1247 -524 1281 452
rect 1405 -524 1439 452
rect 1563 -524 1597 452
rect 1721 -524 1755 452
<< poly >>
rect -1709 545 -1609 561
rect -1709 511 -1693 545
rect -1625 511 -1609 545
rect -1709 464 -1609 511
rect -1551 545 -1451 561
rect -1551 511 -1535 545
rect -1467 511 -1451 545
rect -1551 464 -1451 511
rect -1393 545 -1293 561
rect -1393 511 -1377 545
rect -1309 511 -1293 545
rect -1393 464 -1293 511
rect -1235 545 -1135 561
rect -1235 511 -1219 545
rect -1151 511 -1135 545
rect -1235 464 -1135 511
rect -1077 545 -977 561
rect -1077 511 -1061 545
rect -993 511 -977 545
rect -1077 464 -977 511
rect -919 545 -819 561
rect -919 511 -903 545
rect -835 511 -819 545
rect -919 464 -819 511
rect -761 545 -661 561
rect -761 511 -745 545
rect -677 511 -661 545
rect -761 464 -661 511
rect -603 545 -503 561
rect -603 511 -587 545
rect -519 511 -503 545
rect -603 464 -503 511
rect -445 545 -345 561
rect -445 511 -429 545
rect -361 511 -345 545
rect -445 464 -345 511
rect -287 545 -187 561
rect -287 511 -271 545
rect -203 511 -187 545
rect -287 464 -187 511
rect -129 545 -29 561
rect -129 511 -113 545
rect -45 511 -29 545
rect -129 464 -29 511
rect 29 545 129 561
rect 29 511 45 545
rect 113 511 129 545
rect 29 464 129 511
rect 187 545 287 561
rect 187 511 203 545
rect 271 511 287 545
rect 187 464 287 511
rect 345 545 445 561
rect 345 511 361 545
rect 429 511 445 545
rect 345 464 445 511
rect 503 545 603 561
rect 503 511 519 545
rect 587 511 603 545
rect 503 464 603 511
rect 661 545 761 561
rect 661 511 677 545
rect 745 511 761 545
rect 661 464 761 511
rect 819 545 919 561
rect 819 511 835 545
rect 903 511 919 545
rect 819 464 919 511
rect 977 545 1077 561
rect 977 511 993 545
rect 1061 511 1077 545
rect 977 464 1077 511
rect 1135 545 1235 561
rect 1135 511 1151 545
rect 1219 511 1235 545
rect 1135 464 1235 511
rect 1293 545 1393 561
rect 1293 511 1309 545
rect 1377 511 1393 545
rect 1293 464 1393 511
rect 1451 545 1551 561
rect 1451 511 1467 545
rect 1535 511 1551 545
rect 1451 464 1551 511
rect 1609 545 1709 561
rect 1609 511 1625 545
rect 1693 511 1709 545
rect 1609 464 1709 511
rect -1709 -562 -1609 -536
rect -1551 -562 -1451 -536
rect -1393 -562 -1293 -536
rect -1235 -562 -1135 -536
rect -1077 -562 -977 -536
rect -919 -562 -819 -536
rect -761 -562 -661 -536
rect -603 -562 -503 -536
rect -445 -562 -345 -536
rect -287 -562 -187 -536
rect -129 -562 -29 -536
rect 29 -562 129 -536
rect 187 -562 287 -536
rect 345 -562 445 -536
rect 503 -562 603 -536
rect 661 -562 761 -536
rect 819 -562 919 -536
rect 977 -562 1077 -536
rect 1135 -562 1235 -536
rect 1293 -562 1393 -536
rect 1451 -562 1551 -536
rect 1609 -562 1709 -536
<< polycont >>
rect -1693 511 -1625 545
rect -1535 511 -1467 545
rect -1377 511 -1309 545
rect -1219 511 -1151 545
rect -1061 511 -993 545
rect -903 511 -835 545
rect -745 511 -677 545
rect -587 511 -519 545
rect -429 511 -361 545
rect -271 511 -203 545
rect -113 511 -45 545
rect 45 511 113 545
rect 203 511 271 545
rect 361 511 429 545
rect 519 511 587 545
rect 677 511 745 545
rect 835 511 903 545
rect 993 511 1061 545
rect 1151 511 1219 545
rect 1309 511 1377 545
rect 1467 511 1535 545
rect 1625 511 1693 545
<< locali >>
rect -1709 511 -1693 545
rect -1625 511 -1609 545
rect -1551 511 -1535 545
rect -1467 511 -1451 545
rect -1393 511 -1377 545
rect -1309 511 -1293 545
rect -1235 511 -1219 545
rect -1151 511 -1135 545
rect -1077 511 -1061 545
rect -993 511 -977 545
rect -919 511 -903 545
rect -835 511 -819 545
rect -761 511 -745 545
rect -677 511 -661 545
rect -603 511 -587 545
rect -519 511 -503 545
rect -445 511 -429 545
rect -361 511 -345 545
rect -287 511 -271 545
rect -203 511 -187 545
rect -129 511 -113 545
rect -45 511 -29 545
rect 29 511 45 545
rect 113 511 129 545
rect 187 511 203 545
rect 271 511 287 545
rect 345 511 361 545
rect 429 511 445 545
rect 503 511 519 545
rect 587 511 603 545
rect 661 511 677 545
rect 745 511 761 545
rect 819 511 835 545
rect 903 511 919 545
rect 977 511 993 545
rect 1061 511 1077 545
rect 1135 511 1151 545
rect 1219 511 1235 545
rect 1293 511 1309 545
rect 1377 511 1393 545
rect 1451 511 1467 545
rect 1535 511 1551 545
rect 1609 511 1625 545
rect 1693 511 1709 545
rect -1755 452 -1721 468
rect -1755 -540 -1721 -524
rect -1597 452 -1563 468
rect -1597 -540 -1563 -524
rect -1439 452 -1405 468
rect -1439 -540 -1405 -524
rect -1281 452 -1247 468
rect -1281 -540 -1247 -524
rect -1123 452 -1089 468
rect -1123 -540 -1089 -524
rect -965 452 -931 468
rect -965 -540 -931 -524
rect -807 452 -773 468
rect -807 -540 -773 -524
rect -649 452 -615 468
rect -649 -540 -615 -524
rect -491 452 -457 468
rect -491 -540 -457 -524
rect -333 452 -299 468
rect -333 -540 -299 -524
rect -175 452 -141 468
rect -175 -540 -141 -524
rect -17 452 17 468
rect -17 -540 17 -524
rect 141 452 175 468
rect 141 -540 175 -524
rect 299 452 333 468
rect 299 -540 333 -524
rect 457 452 491 468
rect 457 -540 491 -524
rect 615 452 649 468
rect 615 -540 649 -524
rect 773 452 807 468
rect 773 -540 807 -524
rect 931 452 965 468
rect 931 -540 965 -524
rect 1089 452 1123 468
rect 1089 -540 1123 -524
rect 1247 452 1281 468
rect 1247 -540 1281 -524
rect 1405 452 1439 468
rect 1405 -540 1439 -524
rect 1563 452 1597 468
rect 1563 -540 1597 -524
rect 1721 452 1755 468
rect 1721 -540 1755 -524
<< viali >>
rect -1693 511 -1625 545
rect -1535 511 -1467 545
rect -1377 511 -1309 545
rect -1219 511 -1151 545
rect -1061 511 -993 545
rect -903 511 -835 545
rect -745 511 -677 545
rect -587 511 -519 545
rect -429 511 -361 545
rect -271 511 -203 545
rect -113 511 -45 545
rect 45 511 113 545
rect 203 511 271 545
rect 361 511 429 545
rect 519 511 587 545
rect 677 511 745 545
rect 835 511 903 545
rect 993 511 1061 545
rect 1151 511 1219 545
rect 1309 511 1377 545
rect 1467 511 1535 545
rect 1625 511 1693 545
rect -1755 -507 -1721 -214
rect -1597 142 -1563 435
rect -1439 -507 -1405 -214
rect -1281 142 -1247 435
rect -1123 -507 -1089 -214
rect -965 142 -931 435
rect -807 -507 -773 -214
rect -649 142 -615 435
rect -491 -507 -457 -214
rect -333 142 -299 435
rect -175 -507 -141 -214
rect -17 142 17 435
rect 141 -507 175 -214
rect 299 142 333 435
rect 457 -507 491 -214
rect 615 142 649 435
rect 773 -507 807 -214
rect 931 142 965 435
rect 1089 -507 1123 -214
rect 1247 142 1281 435
rect 1405 -507 1439 -214
rect 1563 142 1597 435
rect 1721 -507 1755 -214
<< metal1 >>
rect -1705 545 -1613 551
rect -1705 511 -1693 545
rect -1625 511 -1613 545
rect -1705 505 -1613 511
rect -1547 545 -1455 551
rect -1547 511 -1535 545
rect -1467 511 -1455 545
rect -1547 505 -1455 511
rect -1389 545 -1297 551
rect -1389 511 -1377 545
rect -1309 511 -1297 545
rect -1389 505 -1297 511
rect -1231 545 -1139 551
rect -1231 511 -1219 545
rect -1151 511 -1139 545
rect -1231 505 -1139 511
rect -1073 545 -981 551
rect -1073 511 -1061 545
rect -993 511 -981 545
rect -1073 505 -981 511
rect -915 545 -823 551
rect -915 511 -903 545
rect -835 511 -823 545
rect -915 505 -823 511
rect -757 545 -665 551
rect -757 511 -745 545
rect -677 511 -665 545
rect -757 505 -665 511
rect -599 545 -507 551
rect -599 511 -587 545
rect -519 511 -507 545
rect -599 505 -507 511
rect -441 545 -349 551
rect -441 511 -429 545
rect -361 511 -349 545
rect -441 505 -349 511
rect -283 545 -191 551
rect -283 511 -271 545
rect -203 511 -191 545
rect -283 505 -191 511
rect -125 545 -33 551
rect -125 511 -113 545
rect -45 511 -33 545
rect -125 505 -33 511
rect 33 545 125 551
rect 33 511 45 545
rect 113 511 125 545
rect 33 505 125 511
rect 191 545 283 551
rect 191 511 203 545
rect 271 511 283 545
rect 191 505 283 511
rect 349 545 441 551
rect 349 511 361 545
rect 429 511 441 545
rect 349 505 441 511
rect 507 545 599 551
rect 507 511 519 545
rect 587 511 599 545
rect 507 505 599 511
rect 665 545 757 551
rect 665 511 677 545
rect 745 511 757 545
rect 665 505 757 511
rect 823 545 915 551
rect 823 511 835 545
rect 903 511 915 545
rect 823 505 915 511
rect 981 545 1073 551
rect 981 511 993 545
rect 1061 511 1073 545
rect 981 505 1073 511
rect 1139 545 1231 551
rect 1139 511 1151 545
rect 1219 511 1231 545
rect 1139 505 1231 511
rect 1297 545 1389 551
rect 1297 511 1309 545
rect 1377 511 1389 545
rect 1297 505 1389 511
rect 1455 545 1547 551
rect 1455 511 1467 545
rect 1535 511 1547 545
rect 1455 505 1547 511
rect 1613 545 1705 551
rect 1613 511 1625 545
rect 1693 511 1705 545
rect 1613 505 1705 511
rect -1603 435 -1557 447
rect -1603 142 -1597 435
rect -1563 142 -1557 435
rect -1603 130 -1557 142
rect -1287 435 -1241 447
rect -1287 142 -1281 435
rect -1247 142 -1241 435
rect -1287 130 -1241 142
rect -971 435 -925 447
rect -971 142 -965 435
rect -931 142 -925 435
rect -971 130 -925 142
rect -655 435 -609 447
rect -655 142 -649 435
rect -615 142 -609 435
rect -655 130 -609 142
rect -339 435 -293 447
rect -339 142 -333 435
rect -299 142 -293 435
rect -339 130 -293 142
rect -23 435 23 447
rect -23 142 -17 435
rect 17 142 23 435
rect -23 130 23 142
rect 293 435 339 447
rect 293 142 299 435
rect 333 142 339 435
rect 293 130 339 142
rect 609 435 655 447
rect 609 142 615 435
rect 649 142 655 435
rect 609 130 655 142
rect 925 435 971 447
rect 925 142 931 435
rect 965 142 971 435
rect 925 130 971 142
rect 1241 435 1287 447
rect 1241 142 1247 435
rect 1281 142 1287 435
rect 1241 130 1287 142
rect 1557 435 1603 447
rect 1557 142 1563 435
rect 1597 142 1603 435
rect 1557 130 1603 142
rect -1761 -214 -1715 -202
rect -1761 -507 -1755 -214
rect -1721 -507 -1715 -214
rect -1761 -519 -1715 -507
rect -1445 -214 -1399 -202
rect -1445 -507 -1439 -214
rect -1405 -507 -1399 -214
rect -1445 -519 -1399 -507
rect -1129 -214 -1083 -202
rect -1129 -507 -1123 -214
rect -1089 -507 -1083 -214
rect -1129 -519 -1083 -507
rect -813 -214 -767 -202
rect -813 -507 -807 -214
rect -773 -507 -767 -214
rect -813 -519 -767 -507
rect -497 -214 -451 -202
rect -497 -507 -491 -214
rect -457 -507 -451 -214
rect -497 -519 -451 -507
rect -181 -214 -135 -202
rect -181 -507 -175 -214
rect -141 -507 -135 -214
rect -181 -519 -135 -507
rect 135 -214 181 -202
rect 135 -507 141 -214
rect 175 -507 181 -214
rect 135 -519 181 -507
rect 451 -214 497 -202
rect 451 -507 457 -214
rect 491 -507 497 -214
rect 451 -519 497 -507
rect 767 -214 813 -202
rect 767 -507 773 -214
rect 807 -507 813 -214
rect 767 -519 813 -507
rect 1083 -214 1129 -202
rect 1083 -507 1089 -214
rect 1123 -507 1129 -214
rect 1083 -519 1129 -507
rect 1399 -214 1445 -202
rect 1399 -507 1405 -214
rect 1439 -507 1445 -214
rect 1399 -519 1445 -507
rect 1715 -214 1761 -202
rect 1715 -507 1721 -214
rect 1755 -507 1761 -214
rect 1715 -519 1761 -507
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5 l 0.5 m 1 nf 22 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc -30 viadrn +30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
