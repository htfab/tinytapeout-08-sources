magic
tech sky130A
magscale 1 2
timestamp 1725569918
<< error_p >>
rect -29 481 29 487
rect -29 447 -17 481
rect -29 441 29 447
rect -29 -447 29 -441
rect -29 -481 -17 -447
rect -29 -487 29 -481
<< nwell >>
rect -221 -619 221 619
<< pmos >>
rect -25 -400 25 400
<< pdiff >>
rect -83 388 -25 400
rect -83 -388 -71 388
rect -37 -388 -25 388
rect -83 -400 -25 -388
rect 25 388 83 400
rect 25 -388 37 388
rect 71 -388 83 388
rect 25 -400 83 -388
<< pdiffc >>
rect -71 -388 -37 388
rect 37 -388 71 388
<< nsubdiff >>
rect -185 549 -89 583
rect 89 549 185 583
rect -185 487 -151 549
rect 151 487 185 549
rect -185 -549 -151 -487
rect 151 -549 185 -487
rect -185 -583 -89 -549
rect 89 -583 185 -549
<< nsubdiffcont >>
rect -89 549 89 583
rect -185 -487 -151 487
rect 151 -487 185 487
rect -89 -583 89 -549
<< poly >>
rect -33 481 33 497
rect -33 447 -17 481
rect 17 447 33 481
rect -33 431 33 447
rect -25 400 25 431
rect -25 -431 25 -400
rect -33 -447 33 -431
rect -33 -481 -17 -447
rect 17 -481 33 -447
rect -33 -497 33 -481
<< polycont >>
rect -17 447 17 481
rect -17 -481 17 -447
<< locali >>
rect -185 549 -89 583
rect 89 549 185 583
rect -185 487 -151 549
rect 151 487 185 549
rect -33 447 -17 481
rect 17 447 33 481
rect -71 388 -37 404
rect -71 -404 -37 -388
rect 37 388 71 404
rect 37 -404 71 -388
rect -33 -481 -17 -447
rect 17 -481 33 -447
rect -185 -549 -151 -487
rect 151 -549 185 -487
rect -185 -583 -89 -549
rect 89 -583 185 -549
<< viali >>
rect -17 447 17 481
rect -71 -388 -37 388
rect 37 -388 71 388
rect -17 -481 17 -447
<< metal1 >>
rect -29 481 29 487
rect -29 447 -17 481
rect 17 447 29 481
rect -29 441 29 447
rect -77 388 -31 400
rect -77 -388 -71 388
rect -37 -388 -31 388
rect -77 -400 -31 -388
rect 31 388 77 400
rect 31 -388 37 388
rect 71 -388 77 388
rect 31 -400 77 -388
rect -29 -447 29 -441
rect -29 -481 -17 -447
rect 17 -481 29 -447
rect -29 -487 29 -481
<< properties >>
string FIXED_BBOX -168 -566 168 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
