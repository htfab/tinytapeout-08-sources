* NGSPICE file created from opamp_l_parax.ext - technology: sky130A

.subckt opamp_l_parax VDD VSS in MINUS PLUS opout
X0 opout.t3 a_n2506_n1366.t8 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 VDD.t5 a_n2506_n1366.t0 a_n2506_n1366.t1 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 opout.t4 MINUS.t0 a_n603_n1314# VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=4
X3 a_n2506_n1366.t7 PLUS.t0 a_n603_n1314# VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=4
X4 opout.t5 MINUS.t1 a_n603_n1314# VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=4
X5 a_n603_n1314# in.t2 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X6 a_n2506_n1366.t3 a_n2506_n1366.t2 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X7 a_n603_n1314# PLUS.t1 a_n2506_n1366.t6 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=4
X8 a_n603_n1314# MINUS.t2 opout.t0 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=4
X9 VSS.t1 in.t3 a_n603_n1314# VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X10 a_n603_n1314# PLUS.t2 a_n2506_n1366.t5 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=4
X11 in.t1 in.t0 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X12 VDD.t1 a_n2506_n1366.t9 opout.t2 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X13 a_n603_n1314# MINUS.t3 opout.t1 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=4
X14 a_n2506_n1366.t4 PLUS.t3 a_n603_n1314# VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=4
R0 a_n2506_n1366.n0 a_n2506_n1366.t9 192.738
R1 a_n2506_n1366.n0 a_n2506_n1366.t2 192.602
R2 a_n2506_n1366.n0 a_n2506_n1366.t0 192.475
R3 a_n2506_n1366.n0 a_n2506_n1366.t8 192.475
R4 a_n2506_n1366.n5 a_n2506_n1366.n4 152.282
R5 a_n2506_n1366.n3 a_n2506_n1366.n1 116.352
R6 a_n2506_n1366.n3 a_n2506_n1366.n2 116.275
R7 a_n2506_n1366.n4 a_n2506_n1366.n3 8.96549
R8 a_n2506_n1366.t1 a_n2506_n1366.n5 7.14175
R9 a_n2506_n1366.n5 a_n2506_n1366.t3 7.14175
R10 a_n2506_n1366.n4 a_n2506_n1366.n0 6.8897
R11 a_n2506_n1366.n2 a_n2506_n1366.t6 4.3505
R12 a_n2506_n1366.n2 a_n2506_n1366.t7 4.3505
R13 a_n2506_n1366.n1 a_n2506_n1366.t5 4.3505
R14 a_n2506_n1366.n1 a_n2506_n1366.t4 4.3505
R15 VDD.t0 VDD.n0 269.286
R16 VDD.n5 VDD.t2 257.257
R17 VDD.t6 VDD.t0 174.201
R18 VDD.t4 VDD.t6 174.201
R19 VDD.t2 VDD.t4 174.201
R20 VDD.n4 VDD.t3 159.048
R21 VDD.n1 VDD.t1 159.048
R22 VDD.n3 VDD.n2 151.905
R23 VDD.n2 VDD.t7 7.14175
R24 VDD.n2 VDD.t5 7.14175
R25 VDD VDD.n0 2.00554
R26 VDD VDD.n5 1.85333
R27 VDD.n3 VDD.n1 0.252453
R28 VDD.n4 VDD.n3 0.252453
R29 VDD.n1 VDD.n0 0.0908298
R30 VDD.n5 VDD.n4 0.0791133
R31 opout.n5 opout.n4 164.411
R32 opout.n1 opout.n0 115.919
R33 opout.n3 opout.n2 115.918
R34 opout.n4 opout.t2 7.14175
R35 opout.n4 opout.t3 7.14175
R36 opout opout.n1 6.64164
R37 opout.n5 opout.n3 5.42116
R38 opout.n2 opout.t1 4.3505
R39 opout.n2 opout.t4 4.3505
R40 opout.n0 opout.t0 4.3505
R41 opout.n0 opout.t5 4.3505
R42 opout opout.n5 0.94675
R43 opout.n3 opout.n1 0.819645
R44 MINUS.n0 MINUS.t2 42.596
R45 MINUS.n2 MINUS.t0 42.0779
R46 MINUS.n1 MINUS.t3 42.0779
R47 MINUS.n0 MINUS.t1 42.0779
R48 MINUS.n1 MINUS.n0 0.518616
R49 MINUS.n2 MINUS.n1 0.518616
R50 MINUS MINUS.n2 0.142408
R51 VSS.t7 VSS.t8 1771.56
R52 VSS.t8 VSS.t6 1771.56
R53 VSS.t6 VSS.t9 1771.56
R54 VSS.t9 VSS.t11 1771.56
R55 VSS.t11 VSS.t10 1771.56
R56 VSS.t10 VSS.t12 1771.56
R57 VSS.t12 VSS.t13 1771.56
R58 VSS.n2 VSS.t7 1606.38
R59 VSS.n2 VSS.t2 555.42
R60 VSS.t0 VSS.t4 326.233
R61 VSS.t2 VSS.t0 326.233
R62 VSS VSS.n2 141.355
R63 VSS.n1 VSS.t3 87.1015
R64 VSS.n1 VSS.n0 78.6563
R65 VSS.n0 VSS.t5 8.7005
R66 VSS.n0 VSS.t1 8.7005
R67 VSS VSS.n1 0.0698548
R68 PLUS.n0 PLUS.t2 42.596
R69 PLUS.n2 PLUS.t0 42.0779
R70 PLUS.n1 PLUS.t1 42.0779
R71 PLUS.n0 PLUS.t3 42.0779
R72 PLUS.n1 PLUS.n0 0.518616
R73 PLUS.n2 PLUS.n1 0.518616
R74 PLUS PLUS.n2 0.185283
R75 in.n0 in.t2 284.546
R76 in.n0 in.t3 284.211
R77 in.n1 in.t0 284.211
R78 in.n2 in.t1 87.7302
R79 in.n1 in.n0 0.335246
R80 in in.n1 0.117025
R81 in in.n2 0.116571
R82 in.n2 in 0.0534661
C0 a_n603_n1314# in 0.141878f
C1 PLUS opout 0.19868f
C2 PLUS MINUS 0.117385f
C3 VDD opout 0.369716f
C4 a_n603_n1314# opout 0.600452f
C5 a_n603_n1314# MINUS 1.84219f
C6 VDD PLUS 0.01037f
C7 a_n603_n1314# PLUS 1.81577f
C8 in opout 0.002177f
C9 MINUS in 0.00227f
C10 a_n603_n1314# VDD 0.065088f
C11 MINUS opout 2.48267f
C12 in VSS 1.15051f
C13 MINUS VSS 6.99185f
C14 PLUS VSS 6.552171f
C15 opout VSS 3.947077f
C16 VDD VSS 9.162437f
C17 a_n603_n1314# VSS 3.6882f
C18 PLUS.t2 VSS 0.469811f
C19 PLUS.t3 VSS 0.46642f
C20 PLUS.n0 VSS 0.561543f
C21 PLUS.t1 VSS 0.46642f
C22 PLUS.n1 VSS 0.286086f
C23 PLUS.t0 VSS 0.46642f
C24 PLUS.n2 VSS 0.238019f
C25 MINUS.t2 VSS 0.391505f
C26 MINUS.t1 VSS 0.388648f
C27 MINUS.n0 VSS 0.470428f
C28 MINUS.t3 VSS 0.388648f
C29 MINUS.n1 VSS 0.238384f
C30 MINUS.t0 VSS 0.388648f
C31 MINUS.n2 VSS 0.193179f
C32 opout.t0 VSS 0.017444f
C33 opout.t5 VSS 0.017444f
C34 opout.n0 VSS 0.0585f
C35 opout.n1 VSS 0.416265f
C36 opout.t1 VSS 0.017444f
C37 opout.t4 VSS 0.017444f
C38 opout.n2 VSS 0.0585f
C39 opout.n3 VSS 0.370227f
C40 opout.t2 VSS 0.017444f
C41 opout.t3 VSS 0.017444f
C42 opout.n4 VSS 0.080188f
C43 opout.n5 VSS 1.127f
C44 VDD.n0 VSS 0.36074f
C45 VDD.t1 VSS 0.052394f
C46 VDD.n1 VSS 0.099929f
C47 VDD.t7 VSS 0.010809f
C48 VDD.t5 VSS 0.010809f
C49 VDD.n2 VSS 0.032731f
C50 VDD.n3 VSS 0.137062f
C51 VDD.t3 VSS 0.052394f
C52 VDD.n4 VSS 0.096675f
C53 VDD.t0 VSS 0.433459f
C54 VDD.t6 VSS 0.338256f
C55 VDD.t4 VSS 0.338256f
C56 VDD.t2 VSS 0.388681f
C57 VDD.n5 VSS 0.182558f
C58 a_n2506_n1366.n0 VSS 0.759796f
C59 a_n2506_n1366.t3 VSS 0.030127f
C60 a_n2506_n1366.t9 VSS 0.37312f
C61 a_n2506_n1366.t8 VSS 0.372886f
C62 a_n2506_n1366.t0 VSS 0.372886f
C63 a_n2506_n1366.t2 VSS 0.372985f
C64 a_n2506_n1366.t5 VSS 0.030127f
C65 a_n2506_n1366.t4 VSS 0.030127f
C66 a_n2506_n1366.n1 VSS 0.103906f
C67 a_n2506_n1366.t6 VSS 0.030127f
C68 a_n2506_n1366.t7 VSS 0.030127f
C69 a_n2506_n1366.n2 VSS 0.103275f
C70 a_n2506_n1366.n3 VSS 1.92021f
C71 a_n2506_n1366.n4 VSS 1.24887f
C72 a_n2506_n1366.n5 VSS 0.091295f
C73 a_n2506_n1366.t1 VSS 0.030127f
.ends

