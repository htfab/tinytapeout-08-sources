** sch_path: /home/ttuser/sud_tt08/TT08/xschem/ota5t_1.sch
.subckt ota5t_1 VCC DIFFOUT BIAS MINUS PLUS VSS
*.PININFO PLUS:I MINUS:I VCC:I VSS:I BIAS:I DIFFOUT:O
XM7 DIFFOUT Vleft VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
XM2 Vleft Vleft VCC VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
XM6 Vleft PLUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 m=1
XM4 DIFFOUT MINUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 m=1
XM1 net1 BIAS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=1 m=1
XM3 BIAS BIAS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=1 m=1
XC1 DIFFOUT VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=10
.ends
.end
