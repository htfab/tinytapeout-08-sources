magic
tech sky130A
magscale 1 2
timestamp 1725008763
<< locali >>
rect -150 1129 3430 1150
rect -150 1095 15 1129
rect 49 1095 3430 1129
rect -150 1065 3430 1095
rect -150 959 1016 1065
rect 1122 959 3430 1065
rect -150 880 3430 959
rect 140 720 240 880
rect 360 750 500 760
rect 350 720 530 750
rect 630 720 730 880
rect 1386 574 1432 752
rect 1702 574 1748 752
rect 1790 720 1890 880
rect 2018 574 2064 752
rect -20 500 140 570
rect 728 480 1312 570
rect 349 -154 514 -119
rect 348 -1040 513 -1034
rect 300 -1069 513 -1040
rect 300 -1260 380 -1069
rect 420 -1080 462 -1069
rect 1320 -1200 1380 -960
rect 1000 -1830 1120 -1780
rect -10 -2490 130 -2390
rect 770 -2410 910 -2380
rect 1000 -2410 1040 -1830
rect 1200 -2234 1234 -2072
rect 1516 -2234 1550 -2072
rect 770 -2450 1040 -2410
rect 770 -2480 910 -2450
rect 330 -2730 560 -2690
rect 350 -2790 540 -2730
rect 1590 -2790 1750 -2200
rect 1832 -2234 1866 -2072
rect 2148 -2234 2182 -2072
rect -270 -2948 -164 -2946
rect -50 -2948 2650 -2790
rect -270 -3020 2650 -2948
rect -50 -3110 2650 -3020
<< viali >>
rect 15 1095 49 1129
rect 1016 959 1122 1065
<< metal1 >>
rect -510 1129 260 1150
rect -510 1095 15 1129
rect 49 1095 260 1129
rect -510 1086 260 1095
rect -180 1084 260 1086
rect 918 1065 1206 1148
rect 918 959 1016 1065
rect 1122 959 1206 1065
rect 918 892 1206 959
rect 140 610 730 650
rect 222 607 298 610
rect 250 530 298 607
rect 1548 392 1610 414
rect 1548 340 1551 392
rect 1603 384 1610 392
rect 1603 340 1632 384
rect 1548 328 1632 340
rect 1548 276 1551 328
rect 1603 276 1632 328
rect 1548 264 1632 276
rect 250 200 404 236
rect 154 -258 224 -214
rect 362 -304 404 200
rect 244 -340 404 -304
rect 466 200 618 236
rect 1548 212 1551 264
rect 1603 212 1632 264
rect 1548 200 1632 212
rect 466 -50 508 200
rect 1548 148 1551 200
rect 1603 148 1632 200
rect 1548 136 1632 148
rect 1548 98 1551 136
rect 1550 84 1551 98
rect 1603 84 1632 136
rect 1550 72 1632 84
rect 1550 20 1551 72
rect 1603 20 1632 72
rect 1550 -18 1632 20
rect 1866 373 1924 414
rect 1866 321 1868 373
rect 1920 321 1924 373
rect 1866 309 1924 321
rect 1866 257 1868 309
rect 1920 257 1924 309
rect 1866 245 1924 257
rect 1866 193 1868 245
rect 1920 193 1924 245
rect 1866 181 1924 193
rect 1866 129 1868 181
rect 1920 129 1924 181
rect 1866 117 1924 129
rect 1866 65 1868 117
rect 1920 65 1924 117
rect 1866 53 1924 65
rect 1866 1 1868 53
rect 1920 1 1924 53
rect 1866 -30 1924 1
rect 2182 371 2240 414
rect 2182 319 2184 371
rect 2236 319 2240 371
rect 2182 307 2240 319
rect 2182 255 2184 307
rect 2236 255 2240 307
rect 2182 243 2240 255
rect 2182 191 2184 243
rect 2236 191 2240 243
rect 2182 179 2240 191
rect 2182 127 2184 179
rect 2236 127 2240 179
rect 2182 115 2240 127
rect 2182 63 2184 115
rect 2236 63 2240 115
rect 2182 51 2240 63
rect 2182 -1 2184 51
rect 2236 -1 2240 51
rect 2182 -30 2240 -1
rect 466 -84 1102 -50
rect 466 -302 508 -84
rect 636 -256 720 -214
rect 466 -338 620 -302
rect 1070 -402 1102 -84
rect 1070 -442 2164 -402
rect 1070 -800 1100 -442
rect -34 -882 126 -834
rect 740 -860 890 -812
rect -34 -1034 14 -882
rect 852 -1034 890 -860
rect 1070 -870 1370 -800
rect -34 -1036 890 -1034
rect -34 -1070 888 -1036
rect 580 -1400 640 -1070
rect 950 -1262 1050 -1260
rect 950 -1308 2132 -1262
rect 950 -1310 1050 -1308
rect 250 -2580 290 -2510
rect 150 -2590 740 -2580
rect 950 -2590 990 -1310
rect 1356 -1485 1432 -1464
rect 1674 -1484 1750 -1460
rect 1356 -1537 1357 -1485
rect 1409 -1537 1432 -1485
rect 1356 -1549 1432 -1537
rect 1356 -1601 1357 -1549
rect 1409 -1601 1432 -1549
rect 1356 -1613 1432 -1601
rect 1356 -1665 1357 -1613
rect 1409 -1665 1432 -1613
rect 1356 -1677 1432 -1665
rect 1356 -1729 1357 -1677
rect 1409 -1729 1432 -1677
rect 1356 -1741 1432 -1729
rect 1356 -1793 1357 -1741
rect 1409 -1793 1432 -1741
rect 1356 -1805 1432 -1793
rect 1356 -1857 1357 -1805
rect 1409 -1857 1432 -1805
rect 1356 -1908 1432 -1857
rect 1672 -1487 1750 -1484
rect 1672 -1539 1673 -1487
rect 1725 -1539 1750 -1487
rect 1672 -1551 1750 -1539
rect 1672 -1603 1673 -1551
rect 1725 -1603 1750 -1551
rect 1672 -1615 1750 -1603
rect 1672 -1667 1673 -1615
rect 1725 -1667 1750 -1615
rect 1672 -1679 1750 -1667
rect 1672 -1731 1673 -1679
rect 1725 -1731 1750 -1679
rect 1672 -1743 1750 -1731
rect 1672 -1795 1673 -1743
rect 1725 -1795 1750 -1743
rect 1672 -1807 1750 -1795
rect 1672 -1859 1673 -1807
rect 1725 -1859 1750 -1807
rect 1672 -1862 1750 -1859
rect 1674 -1904 1750 -1862
rect 1990 -1489 2066 -1458
rect 1990 -1541 1991 -1489
rect 2043 -1541 2066 -1489
rect 1990 -1553 2066 -1541
rect 1990 -1605 1991 -1553
rect 2043 -1605 2066 -1553
rect 1990 -1617 2066 -1605
rect 1990 -1669 1991 -1617
rect 2043 -1669 2066 -1617
rect 1990 -1681 2066 -1669
rect 1990 -1733 1991 -1681
rect 2043 -1733 2066 -1681
rect 1990 -1745 2066 -1733
rect 1990 -1797 1991 -1745
rect 2043 -1797 2066 -1745
rect 1990 -1809 2066 -1797
rect 1990 -1861 1991 -1809
rect 2043 -1861 2066 -1809
rect 1990 -1902 2066 -1861
rect 3510 -1880 3590 -790
rect 3510 -1939 10200 -1880
rect 3510 -1991 10134 -1939
rect 10186 -1991 10200 -1939
rect 3510 -2040 10200 -1991
rect 150 -2626 990 -2590
rect -508 -2630 990 -2626
rect -508 -2688 252 -2630
rect -508 -2690 -94 -2688
rect 150 -2690 242 -2688
<< via1 >>
rect 1551 340 1603 392
rect 1551 276 1603 328
rect 1551 212 1603 264
rect 1551 148 1603 200
rect 1551 84 1603 136
rect 1551 20 1603 72
rect 1868 321 1920 373
rect 1868 257 1920 309
rect 1868 193 1920 245
rect 1868 129 1920 181
rect 1868 65 1920 117
rect 1868 1 1920 53
rect 2184 319 2236 371
rect 2184 255 2236 307
rect 2184 191 2236 243
rect 2184 127 2236 179
rect 2184 63 2236 115
rect 2184 -1 2236 51
rect 1357 -1537 1409 -1485
rect 1357 -1601 1409 -1549
rect 1357 -1665 1409 -1613
rect 1357 -1729 1409 -1677
rect 1357 -1793 1409 -1741
rect 1357 -1857 1409 -1805
rect 1673 -1539 1725 -1487
rect 1673 -1603 1725 -1551
rect 1673 -1667 1725 -1615
rect 1673 -1731 1725 -1679
rect 1673 -1795 1725 -1743
rect 1673 -1859 1725 -1807
rect 1991 -1541 2043 -1489
rect 1991 -1605 2043 -1553
rect 1991 -1669 2043 -1617
rect 1991 -1733 2043 -1681
rect 1991 -1797 2043 -1745
rect 1991 -1861 2043 -1809
rect 10134 -1991 10186 -1939
<< metal2 >>
rect 1494 392 2252 414
rect 1494 340 1551 392
rect 1603 373 2252 392
rect 1603 340 1868 373
rect 1494 328 1868 340
rect 1494 276 1551 328
rect 1603 321 1868 328
rect 1920 371 2252 373
rect 1920 321 2184 371
rect 1603 319 2184 321
rect 2236 319 2252 371
rect 1603 309 2252 319
rect 1603 276 1868 309
rect 1494 264 1868 276
rect 1494 212 1551 264
rect 1603 257 1868 264
rect 1920 307 2252 309
rect 1920 257 2184 307
rect 1603 255 2184 257
rect 2236 255 2252 307
rect 1603 245 2252 255
rect 1603 212 1868 245
rect 1494 200 1868 212
rect 1494 148 1551 200
rect 1603 193 1868 200
rect 1920 243 2252 245
rect 1920 193 2184 243
rect 1603 191 2184 193
rect 2236 191 2252 243
rect 1603 181 2252 191
rect 1603 148 1868 181
rect 1494 136 1868 148
rect 1494 84 1551 136
rect 1603 129 1868 136
rect 1920 179 2252 181
rect 1920 129 2184 179
rect 1603 127 2184 129
rect 2236 127 2252 179
rect 1603 117 2252 127
rect 1603 84 1868 117
rect 1494 72 1868 84
rect 1494 20 1551 72
rect 1603 65 1868 72
rect 1920 115 2252 117
rect 1920 65 2184 115
rect 1603 63 2184 65
rect 2236 63 2252 115
rect 1603 53 2252 63
rect 1603 20 1868 53
rect 1494 1 1868 20
rect 1920 51 2252 53
rect 1920 1 2184 51
rect 1494 -1 2184 1
rect 2236 30 2252 51
rect 2236 -1 3240 30
rect 1494 -22 3240 -1
rect 1494 -30 2802 -22
rect 1620 -238 2802 -30
rect 3178 -238 3240 -22
rect 1620 -290 3240 -238
rect 1626 -1442 1956 -290
rect 1284 -1485 2112 -1442
rect 1284 -1537 1357 -1485
rect 1409 -1487 2112 -1485
rect 1409 -1537 1673 -1487
rect 1284 -1539 1673 -1537
rect 1725 -1489 2112 -1487
rect 1725 -1539 1991 -1489
rect 1284 -1541 1991 -1539
rect 2043 -1541 2112 -1489
rect 1284 -1549 2112 -1541
rect 1284 -1601 1357 -1549
rect 1409 -1551 2112 -1549
rect 1409 -1601 1673 -1551
rect 1284 -1603 1673 -1601
rect 1725 -1553 2112 -1551
rect 1725 -1603 1991 -1553
rect 1284 -1605 1991 -1603
rect 2043 -1605 2112 -1553
rect 1284 -1613 2112 -1605
rect 1284 -1665 1357 -1613
rect 1409 -1615 2112 -1613
rect 1409 -1665 1673 -1615
rect 1284 -1667 1673 -1665
rect 1725 -1617 2112 -1615
rect 1725 -1667 1991 -1617
rect 1284 -1669 1991 -1667
rect 2043 -1669 2112 -1617
rect 1284 -1677 2112 -1669
rect 1284 -1729 1357 -1677
rect 1409 -1679 2112 -1677
rect 1409 -1729 1673 -1679
rect 1284 -1731 1673 -1729
rect 1725 -1681 2112 -1679
rect 1725 -1731 1991 -1681
rect 1284 -1733 1991 -1731
rect 2043 -1733 2112 -1681
rect 1284 -1741 2112 -1733
rect 1284 -1793 1357 -1741
rect 1409 -1743 2112 -1741
rect 1409 -1793 1673 -1743
rect 1284 -1795 1673 -1793
rect 1725 -1745 2112 -1743
rect 1725 -1795 1991 -1745
rect 1284 -1797 1991 -1795
rect 2043 -1797 2112 -1745
rect 1284 -1805 2112 -1797
rect 1284 -1857 1357 -1805
rect 1409 -1807 2112 -1805
rect 1409 -1857 1673 -1807
rect 1284 -1859 1673 -1857
rect 1725 -1809 2112 -1807
rect 1725 -1859 1991 -1809
rect 1284 -1861 1991 -1859
rect 2043 -1861 2112 -1809
rect 1284 -1936 2112 -1861
rect 10120 -1937 10200 -1880
rect 10120 -1993 10132 -1937
rect 10188 -1993 10200 -1937
rect 10120 -2040 10200 -1993
<< via2 >>
rect 2802 -238 3178 -22
rect 10132 -1939 10188 -1937
rect 10132 -1991 10134 -1939
rect 10134 -1991 10186 -1939
rect 10186 -1991 10188 -1939
rect 10132 -1993 10188 -1991
<< metal3 >>
rect 2730 -18 3240 30
rect 2730 -242 2798 -18
rect 3182 -242 3240 -18
rect 2730 -290 3240 -242
rect 10120 -1937 10200 -1380
rect 10120 -1993 10132 -1937
rect 10188 -1993 10200 -1937
rect 10120 -2040 10200 -1993
<< via3 >>
rect 2798 -22 3182 -18
rect 2798 -238 2802 -22
rect 2802 -238 3178 -22
rect 3178 -238 3182 -22
rect 2798 -242 3182 -238
<< metal4 >>
rect 2730 -18 4350 30
rect 2730 -242 2798 -18
rect 3182 -242 4350 -18
rect 2730 -290 4350 -242
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
timestamp 1725008763
transform 1 0 7026 0 1 1250
box -3186 -3040 3186 3040
use sky130_fd_pr__nfet_01v8_3374SR  sky130_fd_pr__nfet_01v8_3374SR_0
timestamp 1725008763
transform 1 0 678 0 1 -594
box -236 -500 236 500
use sky130_fd_pr__nfet_01v8_3374SR  sky130_fd_pr__nfet_01v8_3374SR_1
timestamp 1725008763
transform 1 0 187 0 1 -594
box -236 -500 236 500
use sky130_fd_pr__nfet_01v8_P56BSY  sky130_fd_pr__nfet_01v8_P56BSY_0
timestamp 1725008763
transform 1 0 1691 0 1 -1700
box -631 -560 631 560
use sky130_fd_pr__nfet_01v8_TATN2L  sky130_fd_pr__nfet_01v8_TATN2L_0
timestamp 1725008763
transform 1 0 686 0 1 -1981
box -236 -769 236 769
use sky130_fd_pr__nfet_01v8_TATN2L  sky130_fd_pr__nfet_01v8_TATN2L_1
timestamp 1725008763
transform 1 0 196 0 1 -1981
box -236 -769 236 769
use sky130_fd_pr__pfet_01v8_PDYTS5  sky130_fd_pr__pfet_01v8_PDYTS5_0
timestamp 1725008763
transform 1 0 676 0 1 369
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_PDYTS5  sky130_fd_pr__pfet_01v8_PDYTS5_1
timestamp 1725008763
transform 1 0 193 0 1 366
box -246 -419 246 419
use sky130_fd_pr__pfet_01v8_U25TY6  sky130_fd_pr__pfet_01v8_U25TY6_0
timestamp 1725008763
transform 1 0 1804 0 1 104
box -562 -684 562 684
use sky130_fd_pr__res_generic_po_VBMG2T  sky130_fd_pr__res_generic_po_VBMG2T_0
timestamp 1725008763
transform 0 1 2446 -1 0 -831
box -189 -1286 189 1286
use sky130_fd_pr__res_xhigh_po_0p69_AV7KHZ  sky130_fd_pr__res_xhigh_po_0p69_AV7KHZ_0
timestamp 1725008763
transform 1 0 -437 0 1 -764
box -225 -2442 225 2442
<< labels >>
rlabel metal1 s 954 1000 954 1000 4 VDD
rlabel locali s 850 -2992 850 -2992 4 VSS
rlabel metal1 s 186 -242 186 -242 4 INP
rlabel metal1 s 674 -242 674 -242 4 INM
rlabel metal2 s 2560 -144 2560 -144 4 OUT
<< end >>
