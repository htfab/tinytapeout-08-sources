magic
tech sky130A
magscale 1 2
timestamp 1725528477
<< pwell >>
rect -1522 -712 1522 712
<< psubdiff >>
rect -1486 642 1486 676
rect -1486 580 -1452 642
rect 1452 580 1486 642
rect -1486 -642 -1452 -580
rect 1452 -642 1486 -580
rect -1486 -676 1486 -642
<< psubdiffcont >>
rect -1486 -580 -1452 580
rect 1452 -580 1486 580
<< xpolycontact >>
rect -1356 114 -1218 546
rect -1356 -546 -1218 -114
rect -1122 114 -984 546
rect -1122 -546 -984 -114
rect -888 114 -750 546
rect -888 -546 -750 -114
rect -654 114 -516 546
rect -654 -546 -516 -114
rect -420 114 -282 546
rect -420 -546 -282 -114
rect -186 114 -48 546
rect -186 -546 -48 -114
rect 48 114 186 546
rect 48 -546 186 -114
rect 282 114 420 546
rect 282 -546 420 -114
rect 516 114 654 546
rect 516 -546 654 -114
rect 750 114 888 546
rect 750 -546 888 -114
rect 984 114 1122 546
rect 984 -546 1122 -114
rect 1218 114 1356 546
rect 1218 -546 1356 -114
<< xpolyres >>
rect -1356 -114 -1218 114
rect -1122 -114 -984 114
rect -888 -114 -750 114
rect -654 -114 -516 114
rect -420 -114 -282 114
rect -186 -114 -48 114
rect 48 -114 186 114
rect 282 -114 420 114
rect 516 -114 654 114
rect 750 -114 888 114
rect 984 -114 1122 114
rect 1218 -114 1356 114
<< locali >>
rect -1486 642 1486 676
rect -1486 580 -1452 642
rect 1452 580 1486 642
rect -1486 -642 -1452 -580
rect 1452 -642 1486 -580
rect -1486 -676 1486 -642
<< viali >>
rect -1340 131 -1234 528
rect -1106 131 -1000 528
rect -872 131 -766 528
rect -638 131 -532 528
rect -404 131 -298 528
rect -170 131 -64 528
rect 64 131 170 528
rect 298 131 404 528
rect 532 131 638 528
rect 766 131 872 528
rect 1000 131 1106 528
rect 1234 131 1340 528
rect -1340 -528 -1234 -131
rect -1106 -528 -1000 -131
rect -872 -528 -766 -131
rect -638 -528 -532 -131
rect -404 -528 -298 -131
rect -170 -528 -64 -131
rect 64 -528 170 -131
rect 298 -528 404 -131
rect 532 -528 638 -131
rect 766 -528 872 -131
rect 1000 -528 1106 -131
rect 1234 -528 1340 -131
<< metal1 >>
rect -1346 528 -1228 540
rect -1346 131 -1340 528
rect -1234 131 -1228 528
rect -1346 119 -1228 131
rect -1112 528 -994 540
rect -1112 131 -1106 528
rect -1000 131 -994 528
rect -1112 119 -994 131
rect -878 528 -760 540
rect -878 131 -872 528
rect -766 131 -760 528
rect -878 119 -760 131
rect -644 528 -526 540
rect -644 131 -638 528
rect -532 131 -526 528
rect -644 119 -526 131
rect -410 528 -292 540
rect -410 131 -404 528
rect -298 131 -292 528
rect -410 119 -292 131
rect -176 528 -58 540
rect -176 131 -170 528
rect -64 131 -58 528
rect -176 119 -58 131
rect 58 528 176 540
rect 58 131 64 528
rect 170 131 176 528
rect 58 119 176 131
rect 292 528 410 540
rect 292 131 298 528
rect 404 131 410 528
rect 292 119 410 131
rect 526 528 644 540
rect 526 131 532 528
rect 638 131 644 528
rect 526 119 644 131
rect 760 528 878 540
rect 760 131 766 528
rect 872 131 878 528
rect 760 119 878 131
rect 994 528 1112 540
rect 994 131 1000 528
rect 1106 131 1112 528
rect 994 119 1112 131
rect 1228 528 1346 540
rect 1228 131 1234 528
rect 1340 131 1346 528
rect 1228 119 1346 131
rect -1346 -131 -1228 -119
rect -1346 -528 -1340 -131
rect -1234 -528 -1228 -131
rect -1346 -540 -1228 -528
rect -1112 -131 -994 -119
rect -1112 -528 -1106 -131
rect -1000 -528 -994 -131
rect -1112 -540 -994 -528
rect -878 -131 -760 -119
rect -878 -528 -872 -131
rect -766 -528 -760 -131
rect -878 -540 -760 -528
rect -644 -131 -526 -119
rect -644 -528 -638 -131
rect -532 -528 -526 -131
rect -644 -540 -526 -528
rect -410 -131 -292 -119
rect -410 -528 -404 -131
rect -298 -528 -292 -131
rect -410 -540 -292 -528
rect -176 -131 -58 -119
rect -176 -528 -170 -131
rect -64 -528 -58 -131
rect -176 -540 -58 -528
rect 58 -131 176 -119
rect 58 -528 64 -131
rect 170 -528 176 -131
rect 58 -540 176 -528
rect 292 -131 410 -119
rect 292 -528 298 -131
rect 404 -528 410 -131
rect 292 -540 410 -528
rect 526 -131 644 -119
rect 526 -528 532 -131
rect 638 -528 644 -131
rect 526 -540 644 -528
rect 760 -131 878 -119
rect 760 -528 766 -131
rect 872 -528 878 -131
rect 760 -540 878 -528
rect 994 -131 1112 -119
rect 994 -528 1000 -131
rect 1106 -528 1112 -131
rect 994 -540 1112 -528
rect 1228 -131 1346 -119
rect 1228 -528 1234 -131
rect 1340 -528 1346 -131
rect 1228 -540 1346 -528
<< properties >>
string FIXED_BBOX -1469 -659 1469 659
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 1.3 m 1 nx 12 wmin 0.690 lmin 0.50 rho 2000 val 4.313k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
