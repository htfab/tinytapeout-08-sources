** sch_path: /home/ttuser/tt08_um_alexjaeger_ringoscillator/xschem/ringosc.sch
.subckt ringosc VDD OUT VSS
*.PININFO VDD:I VSS:I OUT:O
x1 VDD VSS net7 net1 not1
x2 VDD VSS net1 net2 not1
x3 VDD VSS net2 net3 not1
x4 VDD VSS net3 net4 not1
x5 VDD VSS net4 net5 not1
x6 VDD VSS net5 net6 not1
x7 VDD VSS net6 net7 not1
x8 VDD VSS net7 OUT notbig
.ends

* expanding   symbol:  not1.sym # of pins=4
** sym_path: /home/ttuser/tt08_um_alexjaeger_ringoscillator/xschem/not1.sym
** sch_path: /home/ttuser/tt08_um_alexjaeger_ringoscillator/xschem/not1.sch
.subckt not1 VDD VSS IN OUT
*.PININFO OUT:O IN:I VDD:I VSS:I
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=5 W=3 nf=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=3 nf=1 m=1
.ends


* expanding   symbol:  notbig.sym # of pins=4
** sym_path: /home/ttuser/tt08_um_alexjaeger_ringoscillator/xschem/notbig.sym
** sch_path: /home/ttuser/tt08_um_alexjaeger_ringoscillator/xschem/notbig.sch
.subckt notbig VDD VSS IN OUT
*.PININFO OUT:O IN:I VDD:I VSS:I
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 m=1
.ends

.end
