magic
tech sky130A
magscale 1 2
timestamp 1723807217
<< nwell >>
rect 1207 1767 1294 2109
<< locali >>
rect 1802 -2366 1838 -1630
rect 2482 -2366 2516 -1632
<< viali >>
rect 1084 2138 1356 2172
rect 2656 2118 2974 2160
rect 1292 -2564 1708 -2528
rect 2660 -2590 3068 -2554
<< metal1 >>
rect -500 2466 6706 2692
rect 418 1966 578 2466
rect 1010 2172 1432 2466
rect 1900 2402 2084 2466
rect 1894 2218 1900 2402
rect 2084 2218 2090 2402
rect 1010 2138 1084 2172
rect 1356 2138 1432 2172
rect 1010 2128 1432 2138
rect 2620 2160 3018 2466
rect 2620 2118 2656 2160
rect 2974 2118 3018 2160
rect 2620 2112 3018 2118
rect 1806 2090 2156 2098
rect 1054 2064 2156 2090
rect 1054 2018 3010 2064
rect 1806 2008 3010 2018
rect 2132 2002 3010 2008
rect -500 846 162 1046
rect 418 994 1034 1966
rect 1900 1622 2084 1628
rect 2276 1622 2566 1906
rect 2084 1438 2566 1622
rect 1900 1432 2084 1438
rect 1454 1162 1850 1234
rect 2276 1226 2566 1438
rect 6736 1384 6742 1488
rect 6846 1384 6852 1488
rect 3008 1176 3492 1240
rect 1454 1087 2013 1162
rect 1454 1014 1850 1087
rect -38 724 162 846
rect -38 518 162 524
rect -510 136 -312 200
rect -510 67 1130 136
rect -510 0 -312 67
rect 1061 -296 1130 67
rect 1621 77 1676 83
rect 1621 -70 1676 22
rect 1598 -248 1699 -70
rect 1061 -333 1744 -296
rect 1061 -350 1130 -333
rect 1938 -410 2013 1087
rect 3008 1014 3495 1176
rect 2461 22 2467 77
rect 2522 22 2528 77
rect 2467 -164 2522 22
rect 2412 -264 2580 -164
rect 3397 -193 3495 1014
rect 6742 -176 6846 1384
rect 6724 -193 6846 -176
rect -500 -624 -242 -564
rect 1610 -585 1622 -470
rect 1735 -485 2013 -410
rect 3397 -291 6857 -193
rect 3397 -411 3495 -291
rect 2549 -509 3495 -411
rect 6724 -479 6857 -291
rect 6990 -479 7190 -370
rect 2138 -565 2422 -528
rect -500 -703 1127 -624
rect -500 -764 -242 -703
rect 1048 -1042 1127 -703
rect 1263 -635 1622 -585
rect 1263 -800 1313 -635
rect 1610 -670 1622 -635
rect 2043 -615 2422 -565
rect 6724 -612 7193 -479
rect 2043 -778 2093 -615
rect 2138 -652 2422 -615
rect 2042 -784 2094 -778
rect 1256 -852 1262 -800
rect 1314 -852 1320 -800
rect 2042 -842 2094 -836
rect 3108 -845 3187 -823
rect 2438 -878 3187 -845
rect 3108 -1042 3187 -878
rect 1048 -1121 3187 -1042
rect 3396 -1248 3448 -1242
rect 3396 -1306 3448 -1300
rect 2742 -1328 2926 -1326
rect 1420 -1330 2926 -1328
rect 1390 -1396 2926 -1330
rect 1390 -1546 1556 -1396
rect 1420 -1566 1497 -1546
rect 1022 -1914 1258 -1790
rect 2020 -1842 2088 -1396
rect 2742 -1580 2926 -1396
rect 654 -2150 1258 -1914
rect 1676 -2039 1963 -1842
rect 2160 -2039 2166 -1842
rect 411 -2623 417 -2571
rect 472 -2623 478 -2571
rect 419 -4129 469 -2623
rect 654 -3076 890 -2150
rect 1022 -2190 1258 -2150
rect 2198 -2048 2628 -1710
rect 3397 -1842 3447 -1306
rect 3053 -1981 3492 -1842
rect 1264 -2522 1744 -2514
rect 1264 -2528 1746 -2522
rect 1264 -2564 1292 -2528
rect 1708 -2564 1746 -2528
rect 1264 -3076 1746 -2564
rect 654 -3312 1746 -3076
rect -526 -21204 -326 -21188
rect 421 -21204 468 -4129
rect 1264 -6196 1746 -3312
rect 2198 -3708 2364 -2048
rect 2642 -2554 3114 -2544
rect 2642 -2560 2660 -2554
rect 1252 -6240 1746 -6196
rect 1938 -6038 2364 -3708
rect 2640 -2590 2660 -2560
rect 3068 -2560 3114 -2554
rect 3068 -2590 3116 -2560
rect 1252 -21204 1740 -6240
rect 1938 -8564 2370 -6038
rect 2640 -6220 3116 -2590
rect 1938 -8570 2384 -8564
rect 1944 -11292 2384 -8570
rect 1938 -11312 2384 -11292
rect 1938 -18216 2376 -11312
rect 1938 -21204 2364 -18216
rect 2618 -21204 3132 -6220
rect 5286 -21026 5390 -21020
rect 5390 -21130 5574 -21026
rect 5286 -21136 5390 -21130
rect 5470 -21204 5574 -21130
rect -536 -21370 6642 -21204
rect -526 -21388 -326 -21370
<< via1 >>
rect 1900 2218 2084 2402
rect 1900 1438 2084 1622
rect 6742 1384 6846 1488
rect -38 524 162 724
rect 1621 22 1676 77
rect 2467 22 2522 77
rect 1262 -852 1314 -800
rect 2042 -836 2094 -784
rect 3396 -1300 3448 -1248
rect 1963 -2039 2160 -1842
rect 417 -2623 472 -2571
rect 5286 -21130 5390 -21026
<< metal2 >>
rect 1900 2402 2084 2408
rect 1900 1622 2084 2218
rect 6742 1741 6846 1746
rect 6738 1647 6747 1741
rect 6841 1647 6850 1741
rect 1894 1438 1900 1622
rect 2084 1438 2090 1622
rect 6742 1488 6846 1647
rect 6742 1378 6846 1384
rect -44 524 -38 724
rect 162 524 168 724
rect -38 -1718 162 524
rect 2467 77 2522 83
rect 1259 22 1621 77
rect 1676 22 2467 77
rect 1259 -102 1314 22
rect 2467 16 2522 22
rect 417 -157 1314 -102
rect -36 -3417 161 -1718
rect 417 -2571 472 -157
rect 1262 -800 1314 -794
rect 2036 -836 2042 -784
rect 2094 -836 2100 -784
rect 1262 -858 1314 -852
rect 1263 -1249 1313 -858
rect 2043 -1249 2093 -836
rect 3390 -1249 3396 -1248
rect 1263 -1299 3396 -1249
rect 3390 -1300 3396 -1299
rect 3448 -1300 3454 -1248
rect 417 -2629 472 -2623
rect 1963 -1842 2160 -1836
rect 1963 -3417 2160 -2039
rect -36 -3614 2160 -3417
rect 5021 -21026 5115 -21022
rect 5016 -21031 5286 -21026
rect 5016 -21125 5021 -21031
rect 5115 -21125 5286 -21031
rect 5016 -21130 5286 -21125
rect 5390 -21130 5396 -21026
rect 5021 -21134 5115 -21130
<< via2 >>
rect 6747 1647 6841 1741
rect 5021 -21125 5115 -21031
<< metal3 >>
rect 6742 1955 6846 1956
rect 6737 1853 6743 1955
rect 6845 1853 6851 1955
rect 6742 1741 6846 1853
rect 6742 1647 6747 1741
rect 6841 1647 6846 1741
rect 6742 1642 6846 1647
rect 4764 -21027 5120 -21026
rect 4759 -21129 4765 -21027
rect 4867 -21031 5120 -21027
rect 4867 -21125 5021 -21031
rect 5115 -21125 5120 -21031
rect 4867 -21129 5120 -21125
rect 4764 -21130 5120 -21129
<< via3 >>
rect 6743 1853 6845 1955
rect 4765 -21129 4867 -21027
<< metal4 >>
rect 6044 2084 6846 2188
rect 6742 1955 6846 2084
rect 6742 1853 6743 1955
rect 6845 1853 6846 1955
rect 6742 1852 6846 1853
rect 4764 -21027 4868 -20886
rect 4764 -21129 4765 -21027
rect 4867 -21129 4868 -21027
rect 4764 -21130 4868 -21129
use sky130_fd_pr__cap_mim_m3_1_72JAQ7  XC1
timestamp 1723797800
transform 1 0 4962 0 1 -9412
box -1186 -11600 1186 11600
use sky130_fd_pr__nfet_01v8_AHRV9L  XM1
timestamp 1723797800
transform 1 0 2842 0 1 -2016
box -396 -610 396 610
use sky130_fd_pr__pfet_01v8_lvt_GWNSVV  XM2
timestamp 1723797800
transform 1 0 1250 0 1 1487
box -396 -719 396 719
use sky130_fd_pr__nfet_01v8_AHRV9L  XM3
timestamp 1723797800
transform 1 0 1480 0 1 -1988
box -396 -610 396 610
use sky130_fd_pr__nfet_01v8_lvt_8TEWK3  XM4
timestamp 1723797800
transform 1 0 2484 0 1 -602
box -246 -410 246 410
use sky130_fd_pr__nfet_01v8_lvt_8TEWK3  XM6
timestamp 1723797800
transform -1 0 1672 0 1 -574
box -246 -410 246 410
use sky130_fd_pr__pfet_01v8_lvt_GWNSVV  XM7
timestamp 1723797800
transform 1 0 2806 0 1 1469
box -396 -719 396 719
<< labels >>
flabel metal1 6990 -570 7190 -370 0 FreeSans 256 0 0 0 DIFFOUT
port 1 nsew
flabel metal1 -488 2476 -288 2676 0 FreeSans 256 0 0 0 VCC
port 0 nsew
flabel metal1 -500 -764 -300 -564 0 FreeSans 256 0 0 0 MINUS
port 3 nsew
flabel space -510 0 -310 200 0 FreeSans 256 0 0 0 PLUS
port 4 nsew
flabel metal1 -500 846 -300 1046 0 FreeSans 256 0 0 0 BIAS
port 2 nsew
flabel metal1 -526 -21388 -326 -21188 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 1938 -485 2013 1162 0 FreeSans 320 0 0 0 Vleft
<< end >>
