magic
tech sky130A
magscale 1 2
timestamp 1725314430
<< nwell >>
rect -941 -619 941 619
<< pmoslvt >>
rect -745 -400 -545 400
rect -487 -400 -287 400
rect -229 -400 -29 400
rect 29 -400 229 400
rect 287 -400 487 400
rect 545 -400 745 400
<< pdiff >>
rect -803 388 -745 400
rect -803 -388 -791 388
rect -757 -388 -745 388
rect -803 -400 -745 -388
rect -545 388 -487 400
rect -545 -388 -533 388
rect -499 -388 -487 388
rect -545 -400 -487 -388
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect 487 388 545 400
rect 487 -388 499 388
rect 533 -388 545 388
rect 487 -400 545 -388
rect 745 388 803 400
rect 745 -388 757 388
rect 791 -388 803 388
rect 745 -400 803 -388
<< pdiffc >>
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
<< nsubdiff >>
rect -905 549 -809 583
rect 809 549 905 583
rect -905 487 -871 549
rect 871 487 905 549
rect -905 -549 -871 -487
rect 871 -549 905 -487
rect -905 -583 -809 -549
rect 809 -583 905 -549
<< nsubdiffcont >>
rect -809 549 809 583
rect -905 -487 -871 487
rect 871 -487 905 487
rect -809 -583 809 -549
<< poly >>
rect -745 481 -545 497
rect -745 447 -729 481
rect -561 447 -545 481
rect -745 400 -545 447
rect -487 481 -287 497
rect -487 447 -471 481
rect -303 447 -287 481
rect -487 400 -287 447
rect -229 481 -29 497
rect -229 447 -213 481
rect -45 447 -29 481
rect -229 400 -29 447
rect 29 481 229 497
rect 29 447 45 481
rect 213 447 229 481
rect 29 400 229 447
rect 287 481 487 497
rect 287 447 303 481
rect 471 447 487 481
rect 287 400 487 447
rect 545 481 745 497
rect 545 447 561 481
rect 729 447 745 481
rect 545 400 745 447
rect -745 -447 -545 -400
rect -745 -481 -729 -447
rect -561 -481 -545 -447
rect -745 -497 -545 -481
rect -487 -447 -287 -400
rect -487 -481 -471 -447
rect -303 -481 -287 -447
rect -487 -497 -287 -481
rect -229 -447 -29 -400
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect -229 -497 -29 -481
rect 29 -447 229 -400
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 29 -497 229 -481
rect 287 -447 487 -400
rect 287 -481 303 -447
rect 471 -481 487 -447
rect 287 -497 487 -481
rect 545 -447 745 -400
rect 545 -481 561 -447
rect 729 -481 745 -447
rect 545 -497 745 -481
<< polycont >>
rect -729 447 -561 481
rect -471 447 -303 481
rect -213 447 -45 481
rect 45 447 213 481
rect 303 447 471 481
rect 561 447 729 481
rect -729 -481 -561 -447
rect -471 -481 -303 -447
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect 303 -481 471 -447
rect 561 -481 729 -447
<< locali >>
rect -905 549 -809 583
rect 809 549 905 583
rect -905 487 -871 549
rect 871 487 905 549
rect -745 447 -729 481
rect -561 447 -545 481
rect -487 447 -471 481
rect -303 447 -287 481
rect -229 447 -213 481
rect -45 447 -29 481
rect 29 447 45 481
rect 213 447 229 481
rect 287 447 303 481
rect 471 447 487 481
rect 545 447 561 481
rect 729 447 745 481
rect -791 388 -757 404
rect -791 -404 -757 -388
rect -533 388 -499 404
rect -533 -404 -499 -388
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect 499 388 533 404
rect 499 -404 533 -388
rect 757 388 791 404
rect 757 -404 791 -388
rect -745 -481 -729 -447
rect -561 -481 -545 -447
rect -487 -481 -471 -447
rect -303 -481 -287 -447
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 287 -481 303 -447
rect 471 -481 487 -447
rect 545 -481 561 -447
rect 729 -481 745 -447
rect -905 -549 -871 -487
rect 871 -549 905 -487
rect -905 -583 -809 -549
rect 809 -583 905 -549
<< viali >>
rect -729 447 -561 481
rect -471 447 -303 481
rect -213 447 -45 481
rect 45 447 213 481
rect 303 447 471 481
rect 561 447 729 481
rect -791 138 -757 371
rect -533 -371 -499 -138
rect -275 138 -241 371
rect -17 -371 17 -138
rect 241 138 275 371
rect 499 -371 533 -138
rect 757 138 791 371
rect -729 -481 -561 -447
rect -471 -481 -303 -447
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect 303 -481 471 -447
rect 561 -481 729 -447
<< metal1 >>
rect -741 481 -549 487
rect -741 447 -729 481
rect -561 447 -549 481
rect -741 441 -549 447
rect -483 481 -291 487
rect -483 447 -471 481
rect -303 447 -291 481
rect -483 441 -291 447
rect -225 481 -33 487
rect -225 447 -213 481
rect -45 447 -33 481
rect -225 441 -33 447
rect 33 481 225 487
rect 33 447 45 481
rect 213 447 225 481
rect 33 441 225 447
rect 291 481 483 487
rect 291 447 303 481
rect 471 447 483 481
rect 291 441 483 447
rect 549 481 741 487
rect 549 447 561 481
rect 729 447 741 481
rect 549 441 741 447
rect -797 371 -751 383
rect -797 138 -791 371
rect -757 138 -751 371
rect -797 126 -751 138
rect -281 371 -235 383
rect -281 138 -275 371
rect -241 138 -235 371
rect -281 126 -235 138
rect 235 371 281 383
rect 235 138 241 371
rect 275 138 281 371
rect 235 126 281 138
rect 751 371 797 383
rect 751 138 757 371
rect 791 138 797 371
rect 751 126 797 138
rect -539 -138 -493 -126
rect -539 -371 -533 -138
rect -499 -371 -493 -138
rect -539 -383 -493 -371
rect -23 -138 23 -126
rect -23 -371 -17 -138
rect 17 -371 23 -138
rect -23 -383 23 -371
rect 493 -138 539 -126
rect 493 -371 499 -138
rect 533 -371 539 -138
rect 493 -383 539 -371
rect -741 -447 -549 -441
rect -741 -481 -729 -447
rect -561 -481 -549 -447
rect -741 -487 -549 -481
rect -483 -447 -291 -441
rect -483 -481 -471 -447
rect -303 -481 -291 -447
rect -483 -487 -291 -481
rect -225 -447 -33 -441
rect -225 -481 -213 -447
rect -45 -481 -33 -447
rect -225 -487 -33 -481
rect 33 -447 225 -441
rect 33 -481 45 -447
rect 213 -481 225 -447
rect 33 -487 225 -481
rect 291 -447 483 -441
rect 291 -481 303 -447
rect 471 -481 483 -447
rect 291 -487 483 -481
rect 549 -447 741 -441
rect 549 -481 561 -447
rect 729 -481 741 -447
rect 549 -487 741 -481
<< properties >>
string FIXED_BBOX -888 -566 888 566
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
