magic
tech sky130A
magscale 1 2
timestamp 1724926688
<< pwell >>
rect -1522 -708 1522 708
<< psubdiff >>
rect -1486 638 -1390 672
rect 1390 638 1486 672
rect -1486 576 -1452 638
rect 1452 576 1486 638
rect -1486 -638 -1452 -576
rect 1452 -638 1486 -576
rect -1486 -672 -1390 -638
rect 1390 -672 1486 -638
<< psubdiffcont >>
rect -1390 638 1390 672
rect -1486 -576 -1452 576
rect 1452 -576 1486 576
rect -1390 -672 1390 -638
<< xpolycontact >>
rect -1356 110 -1218 542
rect -1356 -542 -1218 -110
rect -1122 110 -984 542
rect -1122 -542 -984 -110
rect -888 110 -750 542
rect -888 -542 -750 -110
rect -654 110 -516 542
rect -654 -542 -516 -110
rect -420 110 -282 542
rect -420 -542 -282 -110
rect -186 110 -48 542
rect -186 -542 -48 -110
rect 48 110 186 542
rect 48 -542 186 -110
rect 282 110 420 542
rect 282 -542 420 -110
rect 516 110 654 542
rect 516 -542 654 -110
rect 750 110 888 542
rect 750 -542 888 -110
rect 984 110 1122 542
rect 984 -542 1122 -110
rect 1218 110 1356 542
rect 1218 -542 1356 -110
<< xpolyres >>
rect -1356 -110 -1218 110
rect -1122 -110 -984 110
rect -888 -110 -750 110
rect -654 -110 -516 110
rect -420 -110 -282 110
rect -186 -110 -48 110
rect 48 -110 186 110
rect 282 -110 420 110
rect 516 -110 654 110
rect 750 -110 888 110
rect 984 -110 1122 110
rect 1218 -110 1356 110
<< locali >>
rect -1486 638 -1390 672
rect 1390 638 1486 672
rect -1486 576 -1452 638
rect 1452 576 1486 638
rect -1486 -638 -1452 -576
rect 1452 -638 1486 -576
rect -1486 -672 -1390 -638
rect 1390 -672 1486 -638
<< viali >>
rect -1340 127 -1234 524
rect -1106 127 -1000 524
rect -872 127 -766 524
rect -638 127 -532 524
rect -404 127 -298 524
rect -170 127 -64 524
rect 64 127 170 524
rect 298 127 404 524
rect 532 127 638 524
rect 766 127 872 524
rect 1000 127 1106 524
rect 1234 127 1340 524
rect -1340 -524 -1234 -127
rect -1106 -524 -1000 -127
rect -872 -524 -766 -127
rect -638 -524 -532 -127
rect -404 -524 -298 -127
rect -170 -524 -64 -127
rect 64 -524 170 -127
rect 298 -524 404 -127
rect 532 -524 638 -127
rect 766 -524 872 -127
rect 1000 -524 1106 -127
rect 1234 -524 1340 -127
<< metal1 >>
rect -1346 524 -1228 536
rect -1346 127 -1340 524
rect -1234 127 -1228 524
rect -1346 115 -1228 127
rect -1112 524 -994 536
rect -1112 127 -1106 524
rect -1000 127 -994 524
rect -1112 115 -994 127
rect -878 524 -760 536
rect -878 127 -872 524
rect -766 127 -760 524
rect -878 115 -760 127
rect -644 524 -526 536
rect -644 127 -638 524
rect -532 127 -526 524
rect -644 115 -526 127
rect -410 524 -292 536
rect -410 127 -404 524
rect -298 127 -292 524
rect -410 115 -292 127
rect -176 524 -58 536
rect -176 127 -170 524
rect -64 127 -58 524
rect -176 115 -58 127
rect 58 524 176 536
rect 58 127 64 524
rect 170 127 176 524
rect 58 115 176 127
rect 292 524 410 536
rect 292 127 298 524
rect 404 127 410 524
rect 292 115 410 127
rect 526 524 644 536
rect 526 127 532 524
rect 638 127 644 524
rect 526 115 644 127
rect 760 524 878 536
rect 760 127 766 524
rect 872 127 878 524
rect 760 115 878 127
rect 994 524 1112 536
rect 994 127 1000 524
rect 1106 127 1112 524
rect 994 115 1112 127
rect 1228 524 1346 536
rect 1228 127 1234 524
rect 1340 127 1346 524
rect 1228 115 1346 127
rect -1346 -127 -1228 -115
rect -1346 -524 -1340 -127
rect -1234 -524 -1228 -127
rect -1346 -536 -1228 -524
rect -1112 -127 -994 -115
rect -1112 -524 -1106 -127
rect -1000 -524 -994 -127
rect -1112 -536 -994 -524
rect -878 -127 -760 -115
rect -878 -524 -872 -127
rect -766 -524 -760 -127
rect -878 -536 -760 -524
rect -644 -127 -526 -115
rect -644 -524 -638 -127
rect -532 -524 -526 -127
rect -644 -536 -526 -524
rect -410 -127 -292 -115
rect -410 -524 -404 -127
rect -298 -524 -292 -127
rect -410 -536 -292 -524
rect -176 -127 -58 -115
rect -176 -524 -170 -127
rect -64 -524 -58 -127
rect -176 -536 -58 -524
rect 58 -127 176 -115
rect 58 -524 64 -127
rect 170 -524 176 -127
rect 58 -536 176 -524
rect 292 -127 410 -115
rect 292 -524 298 -127
rect 404 -524 410 -127
rect 292 -536 410 -524
rect 526 -127 644 -115
rect 526 -524 532 -127
rect 638 -524 644 -127
rect 526 -536 644 -524
rect 760 -127 878 -115
rect 760 -524 766 -127
rect 872 -524 878 -127
rect 760 -536 878 -524
rect 994 -127 1112 -115
rect 994 -524 1000 -127
rect 1106 -524 1112 -127
rect 994 -536 1112 -524
rect 1228 -127 1346 -115
rect 1228 -524 1234 -127
rect 1340 -524 1346 -127
rect 1228 -536 1346 -524
<< properties >>
string FIXED_BBOX -1469 -655 1469 655
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 1.26 m 1 nx 12 wmin 0.690 lmin 0.50 rho 2000 val 4.197k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
