magic
tech sky130A
timestamp 1725445236
<< metal1 >>
rect 0 595 100 695
rect 0 290 100 390
rect 640 290 740 390
rect 0 -5 100 95
use vco_inverter  vco_inverter_0
timestamp 1725442979
transform 1 0 -315 0 1 470
box 315 -475 685 225
use vco_inverter  vco_inverter_1
timestamp 1725442979
transform 1 0 55 0 1 470
box 315 -475 685 225
<< labels >>
rlabel metal1 0 645 0 645 7 VDD
port 1 w
rlabel metal1 0 340 0 340 7 Vin
port 3 w
rlabel metal1 0 45 0 45 7 VSS
port 2 w
rlabel metal1 740 340 740 340 3 Vout
port 4 e
<< end >>
