magic
tech sky130A
magscale 1 2
timestamp 1725256794
<< viali >>
rect 19684 1460 22372 1774
<< metal1 >>
rect 26592 13360 30168 13558
rect 30158 13342 30168 13360
rect 30540 13342 30550 13558
rect 194 8658 204 9638
rect 586 8792 596 9638
rect 192 7474 202 8658
rect 586 8476 20964 8792
rect 586 8454 596 8476
rect 584 8110 594 8454
rect 584 7646 4292 8110
rect 584 7474 594 7646
rect 20648 5448 20964 8476
rect 1910 5016 1920 5288
rect 2192 5016 2644 5288
rect 19808 4304 19818 4388
rect 19996 4304 20006 4388
rect 20304 4304 20314 4396
rect 20496 4304 20506 4396
rect 2390 4176 2722 4228
rect 2390 4170 2744 4176
rect 2386 3854 2396 4170
rect 2736 3854 2746 4170
rect 2390 3846 2744 3854
rect 796 1218 806 2254
rect 1186 1820 1196 2254
rect 1186 1426 2955 1820
rect 19672 1774 22384 1780
rect 19672 1460 19684 1774
rect 22372 1460 22384 1774
rect 19672 1454 22384 1460
rect 1186 1340 1196 1426
rect 1188 1320 1198 1340
rect 19964 1320 20268 1454
rect 800 1008 810 1218
rect 1188 1016 20268 1320
rect 1188 1008 1198 1016
<< via1 >>
rect 30168 13342 30540 13558
rect 204 8658 586 9638
rect 202 8454 586 8658
rect 202 7474 584 8454
rect 1920 5016 2192 5288
rect 19818 4304 19996 4388
rect 20314 4304 20496 4396
rect 2396 3854 2736 4170
rect 806 1340 1186 2254
rect 806 1218 1188 1340
rect 810 1008 1188 1218
<< metal2 >>
rect 22530 13868 22714 13878
rect 22530 13624 22714 13634
rect 30168 13558 30540 13568
rect 30168 13332 30540 13342
rect 204 9638 586 9648
rect 202 8658 204 8668
rect 584 8444 586 8454
rect 202 7464 584 7474
rect 1920 5288 2192 5298
rect 1920 5006 2192 5016
rect 19818 4388 19996 4398
rect 19818 4294 19996 4304
rect 20314 4396 20496 4406
rect 20314 4294 20496 4304
rect 2396 4170 2736 4180
rect 2396 3844 2736 3854
rect 806 2254 1186 2264
rect 1186 1340 1188 1350
rect 806 1208 810 1218
rect 810 998 1188 1008
<< via2 >>
rect 22530 13634 22714 13868
rect 30168 13342 30540 13558
rect 204 8658 586 9638
rect 202 8454 586 8658
rect 202 7474 584 8454
rect 1920 5016 2192 5288
rect 19818 4304 19996 4388
rect 20314 4304 20496 4396
rect 2396 3854 2736 4170
rect 806 1340 1186 2254
rect 806 1218 1188 1340
rect 810 1008 1188 1218
<< metal3 >>
rect 204 16482 214 17756
rect 578 17258 588 17756
rect 1974 17258 2828 17260
rect 578 17228 2828 17258
rect 578 16984 2260 17228
rect 2800 16984 2828 17228
rect 578 16972 2828 16984
rect 578 16482 588 16972
rect 22520 13868 22724 13873
rect 22520 13634 22530 13868
rect 22714 13634 22724 13868
rect 22520 13629 22724 13634
rect 30158 13558 30550 13563
rect 30158 13342 30168 13558
rect 30540 13342 30550 13558
rect 30158 13337 30550 13342
rect 794 10142 804 11118
rect 1188 10712 1198 11118
rect 1188 10510 19387 10712
rect 1188 10142 1198 10510
rect 194 9638 596 9643
rect 194 8663 204 9638
rect 192 8658 204 8663
rect 192 7474 202 8658
rect 586 8454 596 9638
rect 23138 9052 23148 9294
rect 23414 9052 23424 9294
rect 584 8449 596 8454
rect 584 7474 594 8449
rect 192 7469 594 7474
rect 1910 5288 2202 5293
rect 1910 5016 1920 5288
rect 2192 5016 2202 5288
rect 1910 5011 2202 5016
rect 20304 4396 20506 4401
rect 19808 4388 20006 4393
rect 19808 4304 19818 4388
rect 19996 4304 20006 4388
rect 19808 4299 20006 4304
rect 20304 4304 20314 4396
rect 20496 4304 20506 4396
rect 20304 4299 20506 4304
rect 2386 4170 2746 4175
rect 2386 3854 2396 4170
rect 2736 3854 2746 4170
rect 2386 3849 2746 3854
rect 796 2254 1196 2259
rect 796 1218 806 2254
rect 1186 1345 1196 2254
rect 1186 1340 1198 1345
rect 796 1213 810 1218
rect 800 1008 810 1213
rect 1188 1008 1198 1340
rect 800 1003 1198 1008
rect 2985 824 3163 829
rect 1920 644 1926 824
rect 2106 823 3186 824
rect 2106 645 2985 823
rect 3163 645 3186 823
rect 2106 644 3186 645
rect 2985 639 3163 644
rect 13796 280 13806 486
rect 14390 468 14400 486
rect 15902 468 15912 486
rect 14390 288 15912 468
rect 14390 280 14400 288
rect 15902 280 15912 288
rect 16496 280 16506 486
rect 17630 212 17810 3978
rect 19342 842 20510 846
rect 19342 838 20512 842
rect 19342 828 20308 838
rect 19342 640 19354 828
rect 19548 650 20308 828
rect 20502 650 20512 838
rect 19548 640 20512 650
rect 23158 748 23338 9052
rect 26262 748 26272 766
rect 19344 638 20306 640
rect 23158 568 26272 748
rect 26262 566 26272 568
rect 26690 566 26700 766
rect 17622 196 18012 212
rect 17622 26 17632 196
rect 18028 26 18038 196
rect 17630 20 17810 26
<< via3 >>
rect 214 16482 578 17756
rect 2260 16984 2800 17228
rect 22530 13634 22714 13868
rect 30168 13342 30540 13558
rect 804 10142 1188 11118
rect 204 8658 586 9638
rect 202 8454 586 8658
rect 23148 9052 23414 9294
rect 202 7474 584 8454
rect 1920 5016 2192 5288
rect 19818 4304 19996 4388
rect 20314 4304 20496 4396
rect 2396 3854 2736 4170
rect 806 1340 1186 2254
rect 806 1218 1188 1340
rect 810 1008 1188 1218
rect 1926 644 2106 824
rect 2985 645 3163 823
rect 13806 280 14390 486
rect 15912 280 16496 486
rect 19354 640 19548 828
rect 20308 650 20502 838
rect 26272 566 26690 766
rect 17632 26 18028 196
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 17756 600 44152
rect 200 16482 214 17756
rect 578 16482 600 17756
rect 200 9638 600 16482
rect 200 8658 204 9638
rect 200 7474 202 8658
rect 586 8454 600 9638
rect 584 7474 600 8454
rect 200 1000 600 7474
rect 800 11118 1200 44152
rect 2259 17228 2801 17229
rect 2259 17216 2260 17228
rect 2258 16988 2260 17216
rect 2259 16984 2260 16988
rect 2800 17216 2801 17228
rect 2800 16988 19602 17216
rect 2800 16984 2801 16988
rect 2259 16983 2801 16984
rect 22529 13868 22715 13869
rect 22529 13826 22530 13868
rect 22522 13634 22530 13826
rect 22714 13826 22715 13868
rect 23250 13826 23406 13838
rect 22714 13634 23406 13826
rect 22522 13632 23406 13634
rect 800 10142 804 11118
rect 1188 10142 1200 11118
rect 800 2254 1200 10142
rect 23250 9295 23406 13632
rect 30167 13558 30541 13559
rect 30167 13342 30168 13558
rect 30540 13542 30541 13558
rect 30540 13342 30542 13542
rect 30167 13341 30542 13342
rect 23147 9294 23415 9295
rect 23147 9052 23148 9294
rect 23414 9052 23415 9294
rect 23147 9051 23415 9052
rect 1919 5288 2193 5289
rect 1919 5016 1920 5288
rect 2192 5016 2193 5288
rect 1919 5015 2193 5016
rect 800 1218 806 2254
rect 1186 1340 1200 2254
rect 800 1008 810 1218
rect 1188 1008 1200 1340
rect 800 1000 1200 1008
rect 1926 825 2106 5015
rect 19816 4389 19996 4418
rect 20313 4396 20497 4397
rect 19816 4388 19997 4389
rect 19816 4304 19818 4388
rect 19996 4304 19997 4388
rect 19816 4303 19997 4304
rect 20313 4304 20314 4396
rect 20496 4304 20497 4396
rect 20313 4303 20497 4304
rect 2395 4170 2737 4171
rect 2395 3854 2396 4170
rect 2736 3854 2737 4170
rect 2395 3853 2737 3854
rect 1925 824 2107 825
rect 1925 644 1926 824
rect 2106 644 2107 824
rect 1925 643 2107 644
rect 2458 468 2638 3853
rect 19353 828 19549 829
rect 19353 824 19354 828
rect 2984 823 19354 824
rect 2984 645 2985 823
rect 3163 645 19354 823
rect 2984 644 19354 645
rect 13805 486 14391 487
rect 13805 468 13806 486
rect 2458 288 13806 468
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 288
rect 13805 280 13806 288
rect 14390 280 14391 486
rect 13805 279 14391 280
rect 14906 0 15086 644
rect 19353 640 19354 644
rect 19548 640 19549 828
rect 19353 639 19549 640
rect 15911 486 16497 487
rect 15911 280 15912 486
rect 16496 468 16497 486
rect 19816 468 19996 4303
rect 20314 839 20494 4303
rect 20307 838 20503 839
rect 20307 650 20308 838
rect 20502 650 20503 838
rect 20307 649 20503 650
rect 20314 640 20494 649
rect 16496 288 19996 468
rect 16496 280 16497 288
rect 15911 279 16497 280
rect 17631 200 18003 212
rect 17630 196 18950 200
rect 17630 26 17632 196
rect 18028 26 18950 196
rect 17630 20 18950 26
rect 18770 0 18950 20
rect 22634 0 22814 4504
rect 26271 766 26691 767
rect 26271 566 26272 766
rect 26690 566 26691 766
rect 26271 565 26691 566
rect 26498 0 26678 565
rect 30362 0 30542 13341
use OPAMP  OPAMP_0 ~/design_submissions_tt08/amr_abdelrahman/magic_sept01
timestamp 1725256412
transform 1 0 3808 0 1 7086
box -1418 -5660 14714 1024
use OPAMP_LAYOUT  OPAMP_LAYOUT_0 ~/design_submissions_tt08/majid_sami/Majid_OpAmp/magic
timestamp 1725008763
transform 1 0 19730 0 1 4568
box -662 -3206 10212 4290
use por  por_0 ~/design_submissions_tt08/khalid_alorayir/magic
timestamp 1725172927
transform 1 0 14962 0 1 6268
box 3566 4220 14642 12130
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
