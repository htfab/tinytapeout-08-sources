magic
tech sky130A
magscale 1 2
timestamp 1725467580
<< nwell >>
rect -581 -498 581 464
<< pmoslvt >>
rect -487 -436 -287 364
rect -229 -436 -29 364
rect 29 -436 229 364
rect 287 -436 487 364
<< pdiff >>
rect -545 352 -487 364
rect -545 -424 -533 352
rect -499 -424 -487 352
rect -545 -436 -487 -424
rect -287 352 -229 364
rect -287 -424 -275 352
rect -241 -424 -229 352
rect -287 -436 -229 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 229 352 287 364
rect 229 -424 241 352
rect 275 -424 287 352
rect 229 -436 287 -424
rect 487 352 545 364
rect 487 -424 499 352
rect 533 -424 545 352
rect 487 -436 545 -424
<< pdiffc >>
rect -533 -424 -499 352
rect -275 -424 -241 352
rect -17 -424 17 352
rect 241 -424 275 352
rect 499 -424 533 352
<< poly >>
rect -487 445 -287 461
rect -487 411 -471 445
rect -303 411 -287 445
rect -487 364 -287 411
rect -229 445 -29 461
rect -229 411 -213 445
rect -45 411 -29 445
rect -229 364 -29 411
rect 29 445 229 461
rect 29 411 45 445
rect 213 411 229 445
rect 29 364 229 411
rect 287 445 487 461
rect 287 411 303 445
rect 471 411 487 445
rect 287 364 487 411
rect -487 -462 -287 -436
rect -229 -462 -29 -436
rect 29 -462 229 -436
rect 287 -462 487 -436
<< polycont >>
rect -471 411 -303 445
rect -213 411 -45 445
rect 45 411 213 445
rect 303 411 471 445
<< locali >>
rect -487 411 -471 445
rect -303 411 -287 445
rect -229 411 -213 445
rect -45 411 -29 445
rect 29 411 45 445
rect 213 411 229 445
rect 287 411 303 445
rect 471 411 487 445
rect -533 352 -499 368
rect -533 -440 -499 -424
rect -275 352 -241 368
rect -275 -440 -241 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 241 352 275 368
rect 241 -440 275 -424
rect 499 352 533 368
rect 499 -440 533 -424
<< viali >>
rect -471 411 -303 445
rect -213 411 -45 445
rect 45 411 213 445
rect 303 411 471 445
rect -533 102 -499 335
rect -275 -407 -241 -174
rect -17 102 17 335
rect 241 -407 275 -174
rect 499 102 533 335
<< metal1 >>
rect -483 445 -291 451
rect -483 411 -471 445
rect -303 411 -291 445
rect -483 405 -291 411
rect -225 445 -33 451
rect -225 411 -213 445
rect -45 411 -33 445
rect -225 405 -33 411
rect 33 445 225 451
rect 33 411 45 445
rect 213 411 225 445
rect 33 405 225 411
rect 291 445 483 451
rect 291 411 303 445
rect 471 411 483 445
rect 291 405 483 411
rect -539 335 -493 347
rect -539 102 -533 335
rect -499 102 -493 335
rect -539 90 -493 102
rect -23 335 23 347
rect -23 102 -17 335
rect 17 102 23 335
rect -23 90 23 102
rect 493 335 539 347
rect 493 102 499 335
rect 533 102 539 335
rect 493 90 539 102
rect -281 -174 -235 -162
rect -281 -407 -275 -174
rect -241 -407 -235 -174
rect -281 -419 -235 -407
rect 235 -174 281 -162
rect 235 -407 241 -174
rect 275 -407 281 -174
rect 235 -419 281 -407
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
