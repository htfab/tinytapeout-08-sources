magic
tech sky130A
magscale 1 2
timestamp 1725314430
<< nwell >>
rect -839 -498 839 464
<< pmoslvt >>
rect -745 -436 -545 364
rect -487 -436 -287 364
rect -229 -436 -29 364
rect 29 -436 229 364
rect 287 -436 487 364
rect 545 -436 745 364
<< pdiff >>
rect -803 352 -745 364
rect -803 -424 -791 352
rect -757 -424 -745 352
rect -803 -436 -745 -424
rect -545 352 -487 364
rect -545 -424 -533 352
rect -499 -424 -487 352
rect -545 -436 -487 -424
rect -287 352 -229 364
rect -287 -424 -275 352
rect -241 -424 -229 352
rect -287 -436 -229 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 229 352 287 364
rect 229 -424 241 352
rect 275 -424 287 352
rect 229 -436 287 -424
rect 487 352 545 364
rect 487 -424 499 352
rect 533 -424 545 352
rect 487 -436 545 -424
rect 745 352 803 364
rect 745 -424 757 352
rect 791 -424 803 352
rect 745 -436 803 -424
<< pdiffc >>
rect -791 -424 -757 352
rect -533 -424 -499 352
rect -275 -424 -241 352
rect -17 -424 17 352
rect 241 -424 275 352
rect 499 -424 533 352
rect 757 -424 791 352
<< poly >>
rect -745 445 -545 461
rect -745 411 -729 445
rect -561 411 -545 445
rect -745 364 -545 411
rect -487 445 -287 461
rect -487 411 -471 445
rect -303 411 -287 445
rect -487 364 -287 411
rect -229 445 -29 461
rect -229 411 -213 445
rect -45 411 -29 445
rect -229 364 -29 411
rect 29 445 229 461
rect 29 411 45 445
rect 213 411 229 445
rect 29 364 229 411
rect 287 445 487 461
rect 287 411 303 445
rect 471 411 487 445
rect 287 364 487 411
rect 545 445 745 461
rect 545 411 561 445
rect 729 411 745 445
rect 545 364 745 411
rect -745 -462 -545 -436
rect -487 -462 -287 -436
rect -229 -462 -29 -436
rect 29 -462 229 -436
rect 287 -462 487 -436
rect 545 -462 745 -436
<< polycont >>
rect -729 411 -561 445
rect -471 411 -303 445
rect -213 411 -45 445
rect 45 411 213 445
rect 303 411 471 445
rect 561 411 729 445
<< locali >>
rect -745 411 -729 445
rect -561 411 -545 445
rect -487 411 -471 445
rect -303 411 -287 445
rect -229 411 -213 445
rect -45 411 -29 445
rect 29 411 45 445
rect 213 411 229 445
rect 287 411 303 445
rect 471 411 487 445
rect 545 411 561 445
rect 729 411 745 445
rect -791 352 -757 368
rect -791 -440 -757 -424
rect -533 352 -499 368
rect -533 -440 -499 -424
rect -275 352 -241 368
rect -275 -440 -241 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 241 352 275 368
rect 241 -440 275 -424
rect 499 352 533 368
rect 499 -440 533 -424
rect 757 352 791 368
rect 757 -440 791 -424
<< viali >>
rect -729 411 -561 445
rect -471 411 -303 445
rect -213 411 -45 445
rect 45 411 213 445
rect 303 411 471 445
rect 561 411 729 445
rect -791 102 -757 335
rect -533 -407 -499 -174
rect -275 102 -241 335
rect -17 -407 17 -174
rect 241 102 275 335
rect 499 -407 533 -174
rect 757 102 791 335
<< metal1 >>
rect -741 445 -549 451
rect -741 411 -729 445
rect -561 411 -549 445
rect -741 405 -549 411
rect -483 445 -291 451
rect -483 411 -471 445
rect -303 411 -291 445
rect -483 405 -291 411
rect -225 445 -33 451
rect -225 411 -213 445
rect -45 411 -33 445
rect -225 405 -33 411
rect 33 445 225 451
rect 33 411 45 445
rect 213 411 225 445
rect 33 405 225 411
rect 291 445 483 451
rect 291 411 303 445
rect 471 411 483 445
rect 291 405 483 411
rect 549 445 741 451
rect 549 411 561 445
rect 729 411 741 445
rect 549 405 741 411
rect -797 335 -751 347
rect -797 102 -791 335
rect -757 102 -751 335
rect -797 90 -751 102
rect -281 335 -235 347
rect -281 102 -275 335
rect -241 102 -235 335
rect -281 90 -235 102
rect 235 335 281 347
rect 235 102 241 335
rect 275 102 281 335
rect 235 90 281 102
rect 751 335 797 347
rect 751 102 757 335
rect 791 102 797 335
rect 751 90 797 102
rect -539 -174 -493 -162
rect -539 -407 -533 -174
rect -499 -407 -493 -174
rect -539 -419 -493 -407
rect -23 -174 23 -162
rect -23 -407 -17 -174
rect 17 -407 23 -174
rect -23 -419 23 -407
rect 493 -174 539 -162
rect 493 -407 499 -174
rect 533 -407 539 -174
rect 493 -419 539 -407
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
