magic
tech sky130A
magscale 1 2
timestamp 1725190886
<< pwell >>
rect -1883 -979 1883 979
<< nmoslvt >>
rect -1687 -769 -887 831
rect -829 -769 -29 831
rect 29 -769 829 831
rect 887 -769 1687 831
<< ndiff >>
rect -1745 819 -1687 831
rect -1745 -757 -1733 819
rect -1699 -757 -1687 819
rect -1745 -769 -1687 -757
rect -887 819 -829 831
rect -887 -757 -875 819
rect -841 -757 -829 819
rect -887 -769 -829 -757
rect -29 819 29 831
rect -29 -757 -17 819
rect 17 -757 29 819
rect -29 -769 29 -757
rect 829 819 887 831
rect 829 -757 841 819
rect 875 -757 887 819
rect 829 -769 887 -757
rect 1687 819 1745 831
rect 1687 -757 1699 819
rect 1733 -757 1745 819
rect 1687 -769 1745 -757
<< ndiffc >>
rect -1733 -757 -1699 819
rect -875 -757 -841 819
rect -17 -757 17 819
rect 841 -757 875 819
rect 1699 -757 1733 819
<< psubdiff >>
rect -1847 909 1847 943
rect -1847 847 -1813 909
rect 1813 847 1847 909
rect -1847 -909 -1813 -847
rect 1813 -909 1847 -847
rect -1847 -943 1847 -909
<< psubdiffcont >>
rect -1847 -847 -1813 847
rect 1813 -847 1847 847
<< poly >>
rect -1687 831 -887 857
rect -829 831 -29 857
rect 29 831 829 857
rect 887 831 1687 857
rect -1687 -807 -887 -769
rect -1687 -841 -1671 -807
rect -903 -841 -887 -807
rect -1687 -857 -887 -841
rect -829 -807 -29 -769
rect -829 -841 -813 -807
rect -45 -841 -29 -807
rect -829 -857 -29 -841
rect 29 -807 829 -769
rect 29 -841 45 -807
rect 813 -841 829 -807
rect 29 -857 829 -841
rect 887 -807 1687 -769
rect 887 -841 903 -807
rect 1671 -841 1687 -807
rect 887 -857 1687 -841
<< polycont >>
rect -1671 -841 -903 -807
rect -813 -841 -45 -807
rect 45 -841 813 -807
rect 903 -841 1671 -807
<< locali >>
rect -1847 909 1847 943
rect -1847 847 -1813 909
rect 1813 847 1847 909
rect -1733 819 -1699 835
rect -1733 -773 -1699 -757
rect -875 819 -841 835
rect -875 -773 -841 -757
rect -17 819 17 835
rect -17 -773 17 -757
rect 841 819 875 835
rect 841 -773 875 -757
rect 1699 819 1733 835
rect 1699 -773 1733 -757
rect -1687 -841 -1671 -807
rect -903 -841 -887 -807
rect -829 -841 -813 -807
rect -45 -841 -29 -807
rect 29 -841 45 -807
rect 813 -841 829 -807
rect 887 -841 903 -807
rect 1671 -841 1687 -807
rect -1847 -909 -1813 -847
rect 1813 -909 1847 -847
rect -1847 -943 1847 -909
<< viali >>
rect -1733 -740 -1699 -267
rect -875 329 -841 802
rect -17 -740 17 -267
rect 841 329 875 802
rect 1699 -740 1733 -267
rect -1671 -841 -903 -807
rect -813 -841 -45 -807
rect 45 -841 813 -807
rect 903 -841 1671 -807
<< metal1 >>
rect -881 802 -835 814
rect -881 329 -875 802
rect -841 329 -835 802
rect -881 317 -835 329
rect 835 802 881 814
rect 835 329 841 802
rect 875 329 881 802
rect 835 317 881 329
rect -1739 -267 -1693 -255
rect -1739 -740 -1733 -267
rect -1699 -740 -1693 -267
rect -1739 -752 -1693 -740
rect -23 -267 23 -255
rect -23 -740 -17 -267
rect 17 -740 23 -267
rect -23 -752 23 -740
rect 1693 -267 1739 -255
rect 1693 -740 1699 -267
rect 1733 -740 1739 -267
rect 1693 -752 1739 -740
rect -1683 -807 -891 -801
rect -1683 -841 -1671 -807
rect -903 -841 -891 -807
rect -1683 -847 -891 -841
rect -825 -807 -33 -801
rect -825 -841 -813 -807
rect -45 -841 -33 -807
rect -825 -847 -33 -841
rect 33 -807 825 -801
rect 33 -841 45 -807
rect 813 -841 825 -807
rect 33 -847 825 -841
rect 891 -807 1683 -801
rect 891 -841 903 -807
rect 1671 -841 1683 -807
rect 891 -847 1683 -841
<< properties >>
string FIXED_BBOX -1830 -926 1830 926
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8 l 4 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -30 viadrn +30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
