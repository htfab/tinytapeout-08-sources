** sch_path: /home/ttuser/tt08_bgr/xschem/BGRwOpampRes.sch
**.subckt BGRwOpampRes
XQ1 VSS VSS MINUS sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ2 VSS VSS net5 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=29
XM1 net1 opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vbgr opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V2 VSS GND 0
Vmeas net1 MINUS 0
.save i(vmeas)
Vmeas1 net2 PLUS 0
.save i(vmeas1)
.save v(vdd)
.save v(net1)
.save v(vdd)
.save v(net2)
.save v(vdd)
.save v(vbgr)
XM4 opout MINUS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Gcm1 PLUS Sop VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 opout Gcm1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(opout)
.save v(sop)
.save v(gcm1)
.save v(sop)
XM10 net3 Gcm2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 Gcm2 Gcm2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Gcm1 Gcm1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.save v(vdd)
.save v(gcm1)
.save v(vdd)
.save v(opout)
.save v(net3)
.save v(vss)
.save v(gcm2)
.save v(vss)
Vmeas3 Sop net3 0
.save i(vmeas3)
XM8 net4 opout VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vmeas2 net4 Gcm2 0
.save i(vmeas2)
.save v(vdd)
.save v(net4)
V3 net6 VSS pwl 0 0 1u 0 4u VDD
E5 TEMPERAT VSS VOL=' temper '
.save v(temperat)
VDD net6 VDD 0
.save i(vdd)
.save v(minus)
.save v(plus)
XR19 net5 PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=0.93 mult=1 m=1
XR3 VSS MINUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6 mult=1 m=1
XR4 VSS Vbgr VSS sky130_fd_pr__res_xhigh_po_0p69 L=12.6 mult=1 m=1
XM12 VSS Vbgr opout opout sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XR2 VSS PLUS VSS sky130_fd_pr__res_xhigh_po_0p35 L=6 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt




* this experimental option enables mos model bin
* selection based on W/NF instead of W
* .options wnflag=1 XMU=0.49 METHOD=GEAR ITL4=100 CHGTOL=1e-15 TRTOL=1 RELTOL=0.0001 VNTOL=0.1u
.param ABSVAR=0.03
.param VCCGAUSS=agauss(1.8, 'ABSVAR', 1)
.param VDD=VCCGAUSS
*.param VDD=1.8
** variation marameters:
* .options savecurrents
.control
  setseed 12
  reset
  let run=1
  dowhile run <= 100
    if run > 1
      reset
      set appendwrite
    end
    * save all
    if run % 3 = 1
      set temp=-40
    end
    if run % 3 = 2
      set temp=27
    end
    if run % 3 = 0
      set temp=125
    end
    echo "Run=$&run, Temp=$temp"
    tran 0.2u 50u
    write lineregulation.raw
    let run = run + 1
  end
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
