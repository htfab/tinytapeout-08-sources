** sch_path: /home/ttuser/test0/tt08-bgr/xschem/opamp_l.sch
.subckt opamp_l VDD VSS in MINUS PLUS opout
*.PININFO VDD:I VSS:I in:I MINUS:I PLUS:I opout:B
XM4 opout MINUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 m=1
XM5 net2 PLUS net1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=16 nf=1 m=1
XM6 opout net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
XM10 net1 in VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=4 nf=1 m=1
XM9 in in VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2 nf=1 m=1
XM7 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=8 nf=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
.ends
.end
