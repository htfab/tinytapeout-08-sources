magic
tech sky130A
magscale 1 2
timestamp 1723727136
<< xpolycontact >>
rect 59 22541 129 22973
rect 225 22541 295 22973
rect 28777 22772 28847 23204
<< ppolyres >>
rect 11015 37088 11251 37158
rect 10683 37010 10919 37080
rect 10351 36836 10587 36906
rect 10019 36661 10255 36731
rect 9687 36487 9923 36557
rect 9355 36313 9591 36383
rect 9023 36138 9259 36208
rect 8691 35964 8927 36034
rect 8359 35808 8595 35860
rect 8691 35808 8761 35964
rect 8857 35953 8927 35964
rect 9023 35953 9093 36138
rect 9189 36087 9259 36138
rect 9355 36087 9425 36313
rect 9521 36213 9591 36313
rect 9687 36213 9757 36487
rect 9853 36329 9923 36487
rect 10019 36329 10089 36661
rect 10185 36436 10255 36661
rect 10351 36436 10421 36836
rect 10517 36534 10587 36836
rect 10683 36534 10753 37010
rect 10849 36623 10919 37010
rect 11015 36623 11085 37088
rect 11181 36704 11251 37088
rect 11347 37088 11583 37158
rect 11347 36704 11417 37088
rect 11513 36777 11583 37088
rect 11679 37088 11915 37158
rect 11679 36777 11749 37088
rect 11513 36707 11749 36777
rect 11845 36842 11915 37088
rect 12011 37088 12247 37158
rect 12011 36842 12081 37088
rect 11845 36772 12081 36842
rect 12177 36898 12247 37088
rect 12343 37088 12579 37158
rect 12343 36898 12413 37088
rect 12177 36828 12413 36898
rect 12509 36947 12579 37088
rect 12675 37088 12911 37158
rect 12675 36947 12745 37088
rect 12509 36877 12745 36947
rect 12841 36987 12911 37088
rect 13007 37088 13243 37158
rect 13007 36987 13077 37088
rect 12841 36917 13077 36987
rect 13173 37020 13243 37088
rect 13339 37088 13575 37158
rect 13339 37020 13409 37088
rect 13173 36950 13409 37020
rect 13505 37045 13575 37088
rect 13671 37088 13907 37158
rect 13671 37045 13741 37088
rect 13505 36975 13741 37045
rect 13837 37063 13907 37088
rect 14003 37088 14239 37158
rect 14003 37063 14073 37088
rect 13837 36993 14073 37063
rect 14169 37072 14239 37088
rect 14335 37088 14571 37158
rect 14335 37072 14405 37088
rect 14169 37002 14405 37072
rect 14501 37074 14571 37088
rect 14667 37088 14903 37158
rect 14667 37074 14737 37088
rect 14501 37004 14737 37074
rect 14833 37068 14903 37088
rect 14999 37088 15235 37158
rect 14999 37068 15069 37088
rect 14833 36998 15069 37068
rect 15165 37055 15235 37088
rect 15331 37088 15567 37158
rect 15331 37055 15401 37088
rect 15165 36985 15401 37055
rect 15497 37034 15567 37088
rect 15663 37088 15899 37158
rect 15663 37034 15733 37088
rect 15497 36964 15733 37034
rect 15829 37005 15899 37088
rect 15995 37088 16231 37158
rect 15995 37005 16065 37088
rect 15829 36935 16065 37005
rect 16161 36968 16231 37088
rect 16327 37088 16563 37158
rect 16327 36968 16397 37088
rect 11181 36634 11417 36704
rect 10849 36553 11085 36623
rect 11513 36541 11749 36611
rect 10517 36464 10753 36534
rect 11181 36468 11417 36538
rect 10185 36366 10421 36436
rect 10849 36387 11085 36457
rect 9853 36259 10089 36329
rect 10517 36298 10753 36368
rect 9521 36143 9757 36213
rect 10185 36200 10421 36270
rect 9189 36017 9425 36087
rect 9853 36093 10089 36163
rect 8857 35883 9093 35953
rect 9521 35977 9757 36047
rect 8359 35790 8761 35808
rect 8027 35653 8263 35686
rect 8359 35653 8429 35790
rect 8525 35738 8761 35790
rect 9189 35851 9425 35921
rect 8027 35616 8429 35653
rect 8857 35717 9093 35787
rect 7695 35488 7931 35511
rect 8027 35488 8097 35616
rect 8193 35583 8429 35616
rect 7695 35441 8097 35488
rect 8525 35572 8761 35642
rect 7363 35312 7599 35337
rect 7695 35312 7765 35441
rect 7861 35418 8097 35441
rect 8193 35417 8429 35487
rect 7363 35267 7765 35312
rect 7031 35124 7267 35163
rect 7363 35124 7433 35267
rect 7529 35242 7765 35267
rect 7861 35252 8097 35322
rect 7031 35093 7433 35124
rect 6699 34925 6935 34988
rect 7031 34925 7101 35093
rect 7197 35054 7433 35093
rect 7529 35076 7765 35146
rect 6699 34918 7101 34925
rect 6367 34744 6603 34814
rect 6035 34570 6271 34640
rect 5703 34395 5939 34465
rect 5371 34221 5607 34291
rect 5039 34047 5275 34117
rect 4707 33873 4943 33943
rect 4375 33698 4611 33768
rect 4043 33524 4279 33594
rect 3711 33323 3947 33393
rect 3379 32789 3615 32859
rect 3047 32157 3283 32227
rect 2715 31525 2951 31595
rect 2383 30892 2619 30962
rect 2051 30272 2287 30330
rect 2383 30272 2453 30892
rect 2549 30785 2619 30892
rect 2715 30785 2785 31525
rect 2881 31254 2951 31525
rect 3047 31254 3117 32157
rect 3213 31686 3283 32157
rect 3379 31686 3449 32789
rect 3545 32086 3615 32789
rect 3711 32086 3781 33323
rect 3877 32459 3947 33323
rect 4043 32459 4113 33524
rect 4209 32807 4279 33524
rect 4375 32807 4445 33698
rect 4541 33132 4611 33698
rect 4707 33132 4777 33873
rect 4873 33438 4943 33873
rect 5039 33438 5109 34047
rect 5205 33725 5275 34047
rect 5371 33725 5441 34221
rect 5537 33994 5607 34221
rect 5703 33994 5773 34395
rect 5869 34248 5939 34395
rect 6035 34248 6105 34570
rect 6201 34488 6271 34570
rect 6367 34488 6437 34744
rect 6533 34713 6603 34744
rect 6699 34713 6769 34918
rect 6865 34855 7101 34918
rect 7197 34888 7433 34958
rect 6533 34643 6769 34713
rect 6865 34689 7101 34759
rect 6201 34418 6437 34488
rect 6533 34477 6769 34547
rect 5869 34178 6105 34248
rect 6201 34252 6437 34322
rect 5537 33924 5773 33994
rect 5869 34012 6105 34082
rect 5205 33655 5441 33725
rect 5537 33758 5773 33828
rect 4873 33368 5109 33438
rect 5205 33489 5441 33559
rect 4541 33062 4777 33132
rect 4873 33202 5109 33272
rect 4209 32737 4445 32807
rect 4541 32896 4777 32966
rect 3877 32389 4113 32459
rect 4209 32571 4445 32641
rect 3545 32016 3781 32086
rect 3877 32223 4113 32293
rect 3213 31616 3449 31686
rect 3545 31850 3781 31920
rect 2881 31184 3117 31254
rect 3213 31450 3449 31520
rect 2549 30715 2785 30785
rect 2881 31018 3117 31088
rect 2051 30260 2453 30272
rect 2051 29706 2121 30260
rect 2217 30202 2453 30260
rect 2549 30549 2785 30619
rect 1719 29636 2121 29706
rect 2217 30036 2453 30106
rect 1719 29073 1789 29636
rect 1387 29003 1789 29073
rect 1885 29470 2121 29540
rect 1055 28363 1291 28433
rect 723 27730 959 27800
rect 391 27098 627 27168
rect 59 26466 295 26536
rect 59 22973 129 26466
rect 225 24658 295 26466
rect 391 24658 461 27098
rect 557 26407 627 27098
rect 723 26407 793 27730
rect 889 27491 959 27730
rect 1055 27491 1125 28363
rect 1221 28348 1291 28363
rect 1387 28348 1457 29003
rect 1221 28278 1457 28348
rect 1553 28837 1789 28907
rect 889 27421 1125 27491
rect 1221 28112 1457 28182
rect 557 26337 793 26407
rect 889 27255 1125 27325
rect 225 24588 461 24658
rect 557 26171 793 26241
rect 225 24422 461 24492
rect 225 22973 295 24422
rect 225 18414 295 22541
rect 391 19689 461 24422
rect 557 19689 627 26171
rect 391 19619 627 19689
rect 391 19453 627 19523
rect 391 18414 461 19453
rect 225 18344 461 18414
rect 557 17782 627 19453
rect 723 18400 793 26171
rect 889 18400 959 27255
rect 723 18330 959 18400
rect 723 18164 959 18234
rect 723 17782 793 18164
rect 557 17712 793 17782
rect 889 17149 959 18164
rect 1055 17448 1125 27255
rect 1221 17448 1291 28112
rect 1055 17378 1291 17448
rect 1055 17212 1291 17282
rect 1055 17149 1125 17212
rect 889 17079 1125 17149
rect 1221 16498 1291 17212
rect 1387 16664 1457 28112
rect 1553 16664 1623 28837
rect 1387 16594 1623 16664
rect 1221 16428 1623 16498
rect 1553 15823 1623 16428
rect 1719 15989 1789 28837
rect 1885 15989 1955 29470
rect 1719 15919 1955 15989
rect 1553 15753 1955 15823
rect 1885 15225 1955 15753
rect 2051 15391 2121 29470
rect 2217 15391 2287 30036
rect 2051 15321 2287 15391
rect 1885 15155 2287 15225
rect 2217 14620 2287 15155
rect 2383 14853 2453 30036
rect 2549 14853 2619 30549
rect 2383 14783 2619 14853
rect 2383 14620 2619 14687
rect 2217 14617 2619 14620
rect 2217 14550 2453 14617
rect 2549 13988 2619 14617
rect 2715 14364 2785 30549
rect 2881 14364 2951 31018
rect 2715 14294 2951 14364
rect 2715 14128 2951 14198
rect 2715 13988 2785 14128
rect 2549 13918 2785 13988
rect 2881 13355 2951 14128
rect 3047 13914 3117 31018
rect 3213 13914 3283 31450
rect 3047 13844 3283 13914
rect 3047 13678 3283 13748
rect 3047 13355 3117 13678
rect 2881 13285 3117 13355
rect 3213 12723 3283 13678
rect 3379 13498 3449 31450
rect 3545 13498 3615 31850
rect 3379 13428 3615 13498
rect 3379 13262 3615 13332
rect 3379 12723 3449 13262
rect 3213 12653 3449 12723
rect 3545 12096 3615 13262
rect 3711 13112 3781 31850
rect 3877 13112 3947 32223
rect 3711 13042 3947 13112
rect 3711 12876 3947 12946
rect 3711 12096 3781 12876
rect 3545 12026 3781 12096
rect 3877 11759 3947 12876
rect 4043 12753 4113 32223
rect 4209 12753 4279 32571
rect 4043 12683 4279 12753
rect 4043 12517 4279 12587
rect 4043 11759 4113 12517
rect 3877 11689 4113 11759
rect 4209 11585 4279 12517
rect 4375 12416 4445 32571
rect 4541 12416 4611 32896
rect 4375 12346 4611 12416
rect 4375 12180 4611 12250
rect 4375 11585 4445 12180
rect 4209 11515 4445 11585
rect 4541 11411 4611 12180
rect 4707 12101 4777 32896
rect 4873 12101 4943 33202
rect 4707 12031 4943 12101
rect 4707 11865 4943 11935
rect 4707 11411 4777 11865
rect 4541 11341 4777 11411
rect 4873 11236 4943 11865
rect 5039 11805 5109 33202
rect 5205 11805 5275 33489
rect 5039 11735 5275 11805
rect 5039 11569 5275 11639
rect 5039 11236 5109 11569
rect 4873 11166 5109 11236
rect 5205 11062 5275 11569
rect 5371 11526 5441 33489
rect 5537 11526 5607 33758
rect 5371 11456 5607 11526
rect 5371 11290 5607 11360
rect 5371 11062 5441 11290
rect 5205 10992 5441 11062
rect 5537 10888 5607 11290
rect 5703 11265 5773 33758
rect 5869 11265 5939 34012
rect 5703 11195 5939 11265
rect 5703 11029 5939 11099
rect 5703 10888 5773 11029
rect 5537 10818 5773 10888
rect 5869 10713 5939 11029
rect 6035 11018 6105 34012
rect 6201 11018 6271 34252
rect 6035 10948 6271 11018
rect 6035 10782 6271 10852
rect 6035 10713 6105 10782
rect 5869 10643 6105 10713
rect 6201 10539 6271 10782
rect 6367 10786 6437 34252
rect 6533 10786 6603 34477
rect 6367 10716 6603 10786
rect 6367 10550 6603 10620
rect 6367 10539 6437 10550
rect 6201 10469 6437 10539
rect 6533 10365 6603 10550
rect 6699 10568 6769 34477
rect 6865 10568 6935 34689
rect 6699 10498 6935 10568
rect 6699 10365 6935 10402
rect 6533 10332 6935 10365
rect 6533 10295 6769 10332
rect 6865 10190 6935 10332
rect 7031 10362 7101 34689
rect 7197 10362 7267 34888
rect 7031 10292 7267 10362
rect 7031 10190 7267 10196
rect 6865 10126 7267 10190
rect 6865 10120 7101 10126
rect 7197 10002 7267 10126
rect 7363 10168 7433 34888
rect 7529 10168 7599 35076
rect 7363 10098 7599 10168
rect 7197 9932 7599 10002
rect 7529 9821 7599 9932
rect 7695 9987 7765 35076
rect 7861 9987 7931 35252
rect 7695 9917 7931 9987
rect 7529 9751 7931 9821
rect 7861 9650 7931 9751
rect 8027 9816 8097 35252
rect 8193 9816 8263 35417
rect 8027 9746 8263 9816
rect 8359 9656 8429 35417
rect 8525 9656 8595 35572
rect 7861 9580 8263 9650
rect 8359 9586 8595 9656
rect 8193 9490 8263 9580
rect 8691 9506 8761 35572
rect 8857 9506 8927 35717
rect 8193 9420 8595 9490
rect 8691 9436 8927 9506
rect 8525 9319 8595 9420
rect 9023 9367 9093 35717
rect 9189 9367 9259 35851
rect 8691 9319 8927 9340
rect 8525 9270 8927 9319
rect 9023 9297 9259 9367
rect 8525 9249 8761 9270
rect 8857 9145 8927 9270
rect 9355 9237 9425 35851
rect 9521 9237 9591 35977
rect 9023 9145 9259 9201
rect 9355 9167 9591 9237
rect 8857 9131 9259 9145
rect 8857 9075 9093 9131
rect 9189 8970 9259 9131
rect 9687 9116 9757 35977
rect 9853 9116 9923 36093
rect 9355 9001 9591 9071
rect 9687 9046 9923 9116
rect 9355 8970 9425 9001
rect 9189 8900 9425 8970
rect 9521 8796 9591 9001
rect 10019 9005 10089 36093
rect 10185 9005 10255 36200
rect 9687 8880 9923 8950
rect 10019 8935 10255 9005
rect 9687 8796 9757 8880
rect 9521 8726 9757 8796
rect 9853 8622 9923 8880
rect 10351 8902 10421 36200
rect 10517 8902 10587 36298
rect 10019 8769 10255 8839
rect 10351 8832 10587 8902
rect 10019 8622 10089 8769
rect 9853 8552 10089 8622
rect 10185 8447 10255 8769
rect 10683 8808 10753 36298
rect 10849 8808 10919 36387
rect 10683 8738 10919 8808
rect 10351 8666 10587 8736
rect 10351 8447 10421 8666
rect 10185 8377 10421 8447
rect 10517 8273 10587 8666
rect 11015 8723 11085 36387
rect 11181 8723 11251 36468
rect 11015 8653 11251 8723
rect 11347 8646 11417 36468
rect 11513 8646 11583 36541
rect 10683 8572 10919 8642
rect 11347 8576 11583 8646
rect 11679 8578 11749 36541
rect 11845 36606 12081 36676
rect 11845 8578 11915 36606
rect 10683 8273 10753 8572
rect 10517 8203 10753 8273
rect 10849 8125 10919 8572
rect 11015 8487 11251 8557
rect 11679 8508 11915 8578
rect 12011 8517 12081 36606
rect 12177 36662 12413 36732
rect 12177 8517 12247 36662
rect 11015 8125 11085 8487
rect 10849 8055 11085 8125
rect 11181 8108 11251 8487
rect 11347 8410 11583 8480
rect 12011 8447 12247 8517
rect 12343 8465 12413 36662
rect 12509 36711 12745 36781
rect 12509 8465 12579 36711
rect 11347 8108 11417 8410
rect 11181 8038 11417 8108
rect 11513 8108 11583 8410
rect 11679 8342 11915 8412
rect 12343 8395 12579 8465
rect 12675 8420 12745 36711
rect 12841 36751 13077 36821
rect 12841 8420 12911 36751
rect 11679 8108 11749 8342
rect 11513 8038 11749 8108
rect 11845 8108 11915 8342
rect 12011 8281 12247 8351
rect 12675 8350 12911 8420
rect 13007 8383 13077 36751
rect 13173 36784 13409 36854
rect 13173 8383 13243 36784
rect 13007 8313 13243 8383
rect 13339 8354 13409 36784
rect 13505 36809 13741 36879
rect 13505 8354 13575 36809
rect 12011 8108 12081 8281
rect 11845 8038 12081 8108
rect 12177 8108 12247 8281
rect 12343 8229 12579 8299
rect 13339 8284 13575 8354
rect 13671 8333 13741 36809
rect 13837 36827 14073 36897
rect 13837 8333 13907 36827
rect 13671 8263 13907 8333
rect 14003 8320 14073 36827
rect 14169 36836 14405 36906
rect 14169 8320 14239 36836
rect 12343 8108 12413 8229
rect 12177 8038 12413 8108
rect 12509 8108 12579 8229
rect 12675 8184 12911 8254
rect 14003 8250 14239 8320
rect 14335 8314 14405 36836
rect 14501 36838 14737 36908
rect 14501 8314 14571 36838
rect 14335 8244 14571 8314
rect 14667 8316 14737 36838
rect 14833 36832 15069 36902
rect 16161 36898 16397 36968
rect 16493 36923 16563 37088
rect 16659 37088 16895 37158
rect 16659 36923 16729 37088
rect 14833 8316 14903 36832
rect 14667 8246 14903 8316
rect 14999 8325 15069 36832
rect 15165 36819 15401 36889
rect 15165 8325 15235 36819
rect 14999 8255 15235 8325
rect 15331 8343 15401 36819
rect 15497 36798 15733 36868
rect 16493 36853 16729 36923
rect 16825 36871 16895 37088
rect 16991 37088 17227 37158
rect 16991 36871 17061 37088
rect 15497 8343 15567 36798
rect 15331 8273 15567 8343
rect 15663 8368 15733 36798
rect 15829 36769 16065 36839
rect 15829 8368 15899 36769
rect 15663 8298 15899 8368
rect 15995 8401 16065 36769
rect 16161 36732 16397 36802
rect 16825 36801 17061 36871
rect 17157 36810 17227 37088
rect 17323 37088 17559 37158
rect 17323 36810 17393 37088
rect 16161 8401 16231 36732
rect 15995 8331 16231 8401
rect 16327 8441 16397 36732
rect 16493 36687 16729 36757
rect 17157 36740 17393 36810
rect 17489 36742 17559 37088
rect 17655 37088 17891 37158
rect 17655 36742 17725 37088
rect 16493 8441 16563 36687
rect 16327 8371 16563 8441
rect 16659 8490 16729 36687
rect 16825 36635 17061 36705
rect 17489 36672 17725 36742
rect 17821 36665 17891 37088
rect 17987 37071 18223 37141
rect 17987 36665 18057 37071
rect 16825 8490 16895 36635
rect 16659 8420 16895 8490
rect 16991 8546 17061 36635
rect 17157 36574 17393 36644
rect 17821 36595 18057 36665
rect 18153 36580 18223 37071
rect 18319 36923 18555 36993
rect 18319 36580 18389 36923
rect 17157 8546 17227 36574
rect 16991 8476 17227 8546
rect 17323 8611 17393 36574
rect 17489 36506 17725 36576
rect 18153 36510 18389 36580
rect 17489 8611 17559 36506
rect 17655 8684 17725 36506
rect 17821 36429 18057 36499
rect 17821 8684 17891 36429
rect 17987 8765 18057 36429
rect 18485 36486 18555 36923
rect 18651 36749 18887 36819
rect 18651 36486 18721 36749
rect 18485 36416 18721 36486
rect 18153 36344 18389 36414
rect 18153 8765 18223 36344
rect 18319 8854 18389 36344
rect 18817 36383 18887 36749
rect 18983 36574 19219 36644
rect 18983 36383 19053 36574
rect 18485 36250 18721 36320
rect 18817 36313 19053 36383
rect 18485 8854 18555 36250
rect 18651 8952 18721 36250
rect 19149 36272 19219 36574
rect 19315 36400 19551 36470
rect 19315 36272 19385 36400
rect 18817 36147 19053 36217
rect 19149 36202 19385 36272
rect 18817 8952 18887 36147
rect 18983 9059 19053 36147
rect 19481 36151 19551 36400
rect 19647 36226 19883 36296
rect 19647 36151 19717 36226
rect 19149 36036 19385 36106
rect 19481 36081 19717 36151
rect 19149 9059 19219 36036
rect 19315 9175 19385 36036
rect 19813 36021 19883 36226
rect 19979 36051 20215 36121
rect 19979 36021 20049 36051
rect 19481 35915 19717 35985
rect 19813 35951 20049 36021
rect 19481 9175 19551 35915
rect 19647 9301 19717 35915
rect 20145 35882 20215 36051
rect 20311 35882 20547 35947
rect 20145 35877 20547 35882
rect 19813 35785 20049 35855
rect 20145 35812 20381 35877
rect 19813 9301 19883 35785
rect 19979 9435 20049 35785
rect 20477 35732 20547 35877
rect 20643 35732 20879 35773
rect 20145 35646 20381 35716
rect 20477 35703 20879 35732
rect 20477 35662 20713 35703
rect 20145 9435 20215 35646
rect 20311 9580 20381 35646
rect 20809 35572 20879 35703
rect 20975 35572 21211 35598
rect 20477 35496 20713 35566
rect 20809 35528 21211 35572
rect 20809 35502 21045 35528
rect 20477 9580 20547 35496
rect 20643 9735 20713 35496
rect 20809 35336 21045 35406
rect 20809 9735 20879 35336
rect 20975 9900 21045 35336
rect 21141 35401 21211 35528
rect 21307 35401 21543 35424
rect 21141 35354 21543 35401
rect 21141 35331 21377 35354
rect 21141 35165 21377 35235
rect 21141 9900 21211 35165
rect 21307 10076 21377 35165
rect 21473 35220 21543 35354
rect 21639 35220 21875 35250
rect 21473 35180 21875 35220
rect 21473 35150 21709 35180
rect 21473 34984 21709 35054
rect 21473 10076 21543 34984
rect 21639 10264 21709 34984
rect 21805 35026 21875 35180
rect 21971 35026 22207 35076
rect 21805 35006 22207 35026
rect 21805 34956 22041 35006
rect 21805 34790 22041 34860
rect 21805 10264 21875 34790
rect 21971 10463 22041 34790
rect 22137 34820 22207 35006
rect 22303 34831 22539 34901
rect 22303 34820 22373 34831
rect 22137 34750 22373 34820
rect 22137 34584 22373 34654
rect 22137 10463 22207 34584
rect 22303 10675 22373 34584
rect 22469 34602 22539 34831
rect 22635 34657 22871 34727
rect 22635 34602 22705 34657
rect 22469 34532 22705 34602
rect 22469 34366 22705 34436
rect 22469 10675 22539 34366
rect 22635 10900 22705 34366
rect 22801 34370 22871 34657
rect 22967 34483 23203 34553
rect 22967 34370 23037 34483
rect 22801 34300 23037 34370
rect 22801 34134 23037 34204
rect 22801 10900 22871 34134
rect 22967 11140 23037 34134
rect 23133 34123 23203 34483
rect 23299 34308 23535 34378
rect 23299 34123 23369 34308
rect 23133 34053 23369 34123
rect 23133 33887 23369 33957
rect 23133 11140 23203 33887
rect 23299 11394 23369 33887
rect 23465 33862 23535 34308
rect 23631 34134 23867 34204
rect 23631 33862 23701 34134
rect 23465 33792 23701 33862
rect 23465 33626 23701 33696
rect 23465 11394 23535 33626
rect 23631 11663 23701 33626
rect 23797 33583 23867 34134
rect 23963 33960 24199 34030
rect 23963 33583 24033 33960
rect 23797 33513 24033 33583
rect 23797 33347 24033 33417
rect 23797 11663 23867 33347
rect 23963 11950 24033 33347
rect 24129 33287 24199 33960
rect 24295 33785 24531 33855
rect 24295 33287 24365 33785
rect 24129 33217 24365 33287
rect 24129 33051 24365 33121
rect 24129 11950 24199 33051
rect 24295 12256 24365 33051
rect 24461 32972 24531 33785
rect 24627 33611 24863 33681
rect 24627 32972 24697 33611
rect 24461 32902 24697 32972
rect 24461 32736 24697 32806
rect 24461 12256 24531 32736
rect 24627 12581 24697 32736
rect 24793 32635 24863 33611
rect 24959 33437 25195 33507
rect 24959 32635 25029 33437
rect 24793 32565 25029 32635
rect 24793 32399 25029 32469
rect 24793 12581 24863 32399
rect 24959 12929 25029 32399
rect 25125 32276 25195 33437
rect 25291 33100 25527 33170
rect 25291 32276 25361 33100
rect 25125 32206 25361 32276
rect 25125 32040 25361 32110
rect 25125 12929 25195 32040
rect 25291 13302 25361 32040
rect 25457 31890 25527 33100
rect 25623 32473 25859 32543
rect 25623 31890 25693 32473
rect 25457 31820 25693 31890
rect 25457 31654 25693 31724
rect 25457 13302 25527 31654
rect 25623 13702 25693 31654
rect 25789 31474 25859 32473
rect 25955 31841 26191 31911
rect 25955 31474 26025 31841
rect 25789 31404 26025 31474
rect 25789 31238 26025 31308
rect 25789 13702 25859 31238
rect 25955 14134 26025 31238
rect 26121 31024 26191 31841
rect 26287 31208 26523 31278
rect 26287 31024 26357 31208
rect 26121 30954 26357 31024
rect 26121 30788 26357 30858
rect 26121 14134 26191 30788
rect 26287 14603 26357 30788
rect 26453 30535 26523 31208
rect 26619 30576 26855 30646
rect 26619 30535 26689 30576
rect 26453 30465 26689 30535
rect 26453 30299 26689 30369
rect 26453 14603 26523 30299
rect 26619 15116 26689 30299
rect 26785 29997 26855 30576
rect 26951 29997 27187 30014
rect 26785 29944 27187 29997
rect 26785 29927 27021 29944
rect 26785 29761 27021 29831
rect 26785 15116 26855 29761
rect 26951 15682 27021 29761
rect 27117 29399 27187 29944
rect 27117 29329 27519 29399
rect 27117 29163 27353 29233
rect 27117 15682 27187 29163
rect 27283 16315 27353 29163
rect 27449 28724 27519 29329
rect 27615 28724 27851 28749
rect 27449 28679 27851 28724
rect 27449 28654 27685 28679
rect 27449 28488 27685 28558
rect 27449 16315 27519 28488
rect 27615 17040 27685 28488
rect 27781 27940 27851 28679
rect 27947 28047 28183 28117
rect 27947 27940 28017 28047
rect 27781 27870 28017 27940
rect 27781 27704 28017 27774
rect 27781 17040 27851 27704
rect 27947 17897 28017 27704
rect 28113 26988 28183 28047
rect 28279 27414 28515 27484
rect 28279 26988 28349 27414
rect 28113 26918 28349 26988
rect 28113 26752 28349 26822
rect 28113 17897 28183 26752
rect 28279 18981 28349 26752
rect 28445 25699 28515 27414
rect 28611 26782 28847 26852
rect 28611 25699 28681 26782
rect 28445 25629 28681 25699
rect 28445 25463 28681 25533
rect 28445 18981 28515 25463
rect 28611 20730 28681 25463
rect 28777 23370 28847 26782
rect 28777 23300 29013 23370
rect 28777 20730 28847 22772
rect 28611 20660 28847 20730
rect 28279 18911 28515 18981
rect 28611 20494 28847 20564
rect 27947 17827 28183 17897
rect 28279 18745 28515 18815
rect 27615 16970 27851 17040
rect 27947 17661 28183 17731
rect 27283 16245 27519 16315
rect 27615 16833 27851 16874
rect 27947 16833 28017 17661
rect 28113 17466 28183 17661
rect 28279 17466 28349 18745
rect 28445 18098 28515 18745
rect 28611 18098 28681 20494
rect 28777 18730 28847 20494
rect 28943 18730 29013 23300
rect 28777 18660 29013 18730
rect 28445 18028 28681 18098
rect 28113 17396 28349 17466
rect 27615 16804 28017 16833
rect 27615 16149 27685 16804
rect 27781 16763 28017 16804
rect 26951 15612 27187 15682
rect 27283 16079 27685 16149
rect 27283 15516 27353 16079
rect 26619 15046 26855 15116
rect 26951 15446 27353 15516
rect 26287 14533 26523 14603
rect 26619 14936 26855 14950
rect 26951 14936 27021 15446
rect 26619 14880 27021 14936
rect 25955 14064 26191 14134
rect 26287 14367 26523 14437
rect 25623 13632 25859 13702
rect 25955 13898 26191 13968
rect 25291 13232 25527 13302
rect 25623 13466 25859 13536
rect 24959 12859 25195 12929
rect 25291 13066 25527 13136
rect 24627 12511 24863 12581
rect 24959 12693 25195 12763
rect 24295 12186 24531 12256
rect 24627 12345 24863 12415
rect 23963 11880 24199 11950
rect 24295 12020 24531 12090
rect 23631 11593 23867 11663
rect 23963 11714 24199 11784
rect 23299 11324 23535 11394
rect 23631 11427 23867 11497
rect 22967 11070 23203 11140
rect 23299 11158 23535 11228
rect 22635 10830 22871 10900
rect 22967 10904 23203 10974
rect 22303 10605 22539 10675
rect 22635 10664 22871 10734
rect 21971 10393 22207 10463
rect 22303 10452 22539 10509
rect 22635 10452 22705 10664
rect 22801 10626 22871 10664
rect 22967 10626 23037 10904
rect 23133 10801 23203 10904
rect 23299 10801 23369 11158
rect 23465 10975 23535 11158
rect 23631 10975 23701 11427
rect 23797 11149 23867 11427
rect 23963 11149 24033 11714
rect 24129 11323 24199 11714
rect 24295 11323 24365 12020
rect 24461 11498 24531 12020
rect 24627 11498 24697 12345
rect 24793 11672 24863 12345
rect 24959 11672 25029 12693
rect 25125 11873 25195 12693
rect 25291 11873 25361 13066
rect 25457 12407 25527 13066
rect 25623 12407 25693 13466
rect 25789 13039 25859 13466
rect 25955 13039 26025 13898
rect 26121 13671 26191 13898
rect 26287 13671 26357 14367
rect 26453 14304 26523 14367
rect 26619 14304 26689 14880
rect 26785 14866 27021 14880
rect 26453 14234 26689 14304
rect 26121 13601 26357 13671
rect 25789 12969 26025 13039
rect 25457 12337 25693 12407
rect 25125 11803 25361 11873
rect 24793 11602 25029 11672
rect 24461 11428 24697 11498
rect 24129 11253 24365 11323
rect 23797 11079 24033 11149
rect 23465 10905 23701 10975
rect 23133 10731 23369 10801
rect 22801 10556 23037 10626
rect 22303 10439 22705 10452
rect 21639 10194 21875 10264
rect 21971 10278 22207 10297
rect 22303 10278 22373 10439
rect 22469 10382 22705 10439
rect 21971 10227 22373 10278
rect 21971 10098 22041 10227
rect 22137 10208 22373 10227
rect 21307 10006 21543 10076
rect 21639 10028 22041 10098
rect 21639 9910 21709 10028
rect 20975 9830 21211 9900
rect 21307 9840 21709 9910
rect 20643 9665 20879 9735
rect 21307 9734 21377 9840
rect 20311 9510 20547 9580
rect 20975 9664 21377 9734
rect 20975 9569 21045 9664
rect 19979 9365 20215 9435
rect 20643 9499 21045 9569
rect 20311 9406 20547 9414
rect 20643 9406 20713 9499
rect 19647 9231 19883 9301
rect 20311 9344 20713 9406
rect 19979 9232 20215 9269
rect 20311 9232 20381 9344
rect 20477 9336 20713 9344
rect 19315 9105 19551 9175
rect 19979 9199 20381 9232
rect 18983 8989 19219 9059
rect 19647 9065 19883 9135
rect 18651 8882 18887 8952
rect 19315 8939 19551 9009
rect 18319 8784 18555 8854
rect 18983 8823 19219 8893
rect 17987 8695 18223 8765
rect 18651 8716 18887 8786
rect 17655 8614 17891 8684
rect 18319 8618 18555 8688
rect 17323 8541 17559 8611
rect 17987 8529 18223 8599
rect 17655 8448 17891 8518
rect 12675 8108 12745 8184
rect 12509 8038 12745 8108
rect 12841 8108 12911 8184
rect 13007 8147 13243 8217
rect 13007 8108 13077 8147
rect 12841 8038 13077 8108
rect 13173 8108 13243 8147
rect 13339 8118 13575 8188
rect 13339 8108 13409 8118
rect 13173 8038 13409 8108
rect 13505 8108 13575 8118
rect 13671 8108 13907 8167
rect 14003 8108 14239 8154
rect 14335 8108 14571 8148
rect 14667 8108 14903 8150
rect 14999 8108 15235 8159
rect 15331 8108 15567 8177
rect 15663 8132 15899 8202
rect 15663 8108 15733 8132
rect 13505 8107 15733 8108
rect 13505 8097 15401 8107
rect 13505 8038 13741 8097
rect 13837 8089 15401 8097
rect 13837 8084 15069 8089
rect 13837 8038 14073 8084
rect 14169 8080 15069 8084
rect 14169 8078 14737 8080
rect 14169 8038 14405 8078
rect 14501 8038 14737 8078
rect 14833 8038 15069 8080
rect 15165 8038 15401 8089
rect 15497 8038 15733 8107
rect 15829 8108 15899 8132
rect 15995 8165 16231 8235
rect 15995 8108 16065 8165
rect 15829 8038 16065 8108
rect 16161 8108 16231 8165
rect 16327 8205 16563 8275
rect 16327 8108 16397 8205
rect 16161 8038 16397 8108
rect 16493 8108 16563 8205
rect 16659 8254 16895 8324
rect 16659 8108 16729 8254
rect 16493 8038 16729 8108
rect 16825 8108 16895 8254
rect 16991 8310 17227 8380
rect 16991 8108 17061 8310
rect 16825 8038 17061 8108
rect 17157 8108 17227 8310
rect 17323 8375 17559 8445
rect 17323 8108 17393 8375
rect 17157 8038 17393 8108
rect 17489 8108 17559 8375
rect 17655 8108 17725 8448
rect 17489 8038 17725 8108
rect 17821 8108 17891 8448
rect 17987 8108 18057 8529
rect 18153 8186 18223 8529
rect 18319 8186 18389 8618
rect 18485 8360 18555 8618
rect 18651 8360 18721 8716
rect 18817 8535 18887 8716
rect 18983 8535 19053 8823
rect 19149 8709 19219 8823
rect 19315 8709 19385 8939
rect 19481 8883 19551 8939
rect 19647 8883 19717 9065
rect 19813 9058 19883 9065
rect 19979 9058 20049 9199
rect 20145 9162 20381 9199
rect 19813 8988 20049 9058
rect 19481 8813 19717 8883
rect 19149 8639 19385 8709
rect 18817 8465 19053 8535
rect 18485 8290 18721 8360
rect 18153 8116 18389 8186
rect 17821 8038 18057 8108
<< labels >>
flabel xpolycontact 59 22541 129 22973 0 FreeSans 400 90 0 0 VPWR
port 1 nsew power bidirectional
flabel xpolycontact 28777 22772 28847 23204 0 FreeSans 400 90 0 0 VGND
port 2 nsew ground bidirectional
flabel xpolycontact 225 22541 295 22973 0 FreeSans 400 90 0 0 VOUT
port 3 nsew analog bidirectional
<< end >>
