** sch_path: /home/ttuser/rr08-analog-ringoscillator/xschem/ring1.sch
**.subckt ring1 out
*.opin out
C1 net1 GND 4f m=1
R1 out net1 500 m=1
V1 net3 GND 1.8
V2 net2 GND 0
Vmeas1 VDD net3 0
.save i(vmeas1)
Vmeas2 VSS net2 0
.save i(vmeas2)
x1 VDD net1 VSS ringosc
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.options savecurrents
.control
save all
tran 0.01n 1000n
write ring1.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  ringosc.sym # of pins=3
** sym_path: /home/ttuser/rr08-analog-ringoscillator/xschem/ringosc.sym
** sch_path: /home/ttuser/rr08-analog-ringoscillator/xschem/ringosc.sch
.subckt ringosc VDD OUT VSS
*.ipin VDD
*.ipin VSS
*.opin OUT
x1 VDD VSS net7 net1 not1
x2 VDD VSS net1 net2 not1
x3 VDD VSS net2 net3 not1
x4 VDD VSS net3 net4 not1
x5 VDD VSS net4 net5 not1
x6 VDD VSS net5 net6 not1
x7 VDD VSS net6 net7 not1
x8 VDD VSS net7 OUT notbig
.ends


* expanding   symbol:  not1.sym # of pins=4
** sym_path: /home/ttuser/rr08-analog-ringoscillator/xschem/not1.sym
** sch_path: /home/ttuser/rr08-analog-ringoscillator/xschem/not1.sch
.subckt not1 VDD VSS IN OUT
*.opin OUT
*.ipin IN
*.ipin VDD
*.ipin VSS
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=5 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  notbig.sym # of pins=4
** sym_path: /home/ttuser/rr08-analog-ringoscillator/xschem/notbig.sym
** sch_path: /home/ttuser/rr08-analog-ringoscillator/xschem/notbig.sch
.subckt notbig VDD VSS IN OUT
*.opin OUT
*.ipin IN
*.ipin VDD
*.ipin VSS
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
