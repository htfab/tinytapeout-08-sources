magic
tech sky130A
magscale 1 2
timestamp 1724939774
<< nwell >>
rect -855 -1098 855 1064
<< pmoslvt >>
rect -761 -1036 -661 964
rect -603 -1036 -503 964
rect -445 -1036 -345 964
rect -287 -1036 -187 964
rect -129 -1036 -29 964
rect 29 -1036 129 964
rect 187 -1036 287 964
rect 345 -1036 445 964
rect 503 -1036 603 964
rect 661 -1036 761 964
<< pdiff >>
rect -819 952 -761 964
rect -819 -1024 -807 952
rect -773 -1024 -761 952
rect -819 -1036 -761 -1024
rect -661 952 -603 964
rect -661 -1024 -649 952
rect -615 -1024 -603 952
rect -661 -1036 -603 -1024
rect -503 952 -445 964
rect -503 -1024 -491 952
rect -457 -1024 -445 952
rect -503 -1036 -445 -1024
rect -345 952 -287 964
rect -345 -1024 -333 952
rect -299 -1024 -287 952
rect -345 -1036 -287 -1024
rect -187 952 -129 964
rect -187 -1024 -175 952
rect -141 -1024 -129 952
rect -187 -1036 -129 -1024
rect -29 952 29 964
rect -29 -1024 -17 952
rect 17 -1024 29 952
rect -29 -1036 29 -1024
rect 129 952 187 964
rect 129 -1024 141 952
rect 175 -1024 187 952
rect 129 -1036 187 -1024
rect 287 952 345 964
rect 287 -1024 299 952
rect 333 -1024 345 952
rect 287 -1036 345 -1024
rect 445 952 503 964
rect 445 -1024 457 952
rect 491 -1024 503 952
rect 445 -1036 503 -1024
rect 603 952 661 964
rect 603 -1024 615 952
rect 649 -1024 661 952
rect 603 -1036 661 -1024
rect 761 952 819 964
rect 761 -1024 773 952
rect 807 -1024 819 952
rect 761 -1036 819 -1024
<< pdiffc >>
rect -807 -1024 -773 952
rect -649 -1024 -615 952
rect -491 -1024 -457 952
rect -333 -1024 -299 952
rect -175 -1024 -141 952
rect -17 -1024 17 952
rect 141 -1024 175 952
rect 299 -1024 333 952
rect 457 -1024 491 952
rect 615 -1024 649 952
rect 773 -1024 807 952
<< poly >>
rect -761 1045 -661 1061
rect -761 1011 -745 1045
rect -677 1011 -661 1045
rect -761 964 -661 1011
rect -603 1045 -503 1061
rect -603 1011 -587 1045
rect -519 1011 -503 1045
rect -603 964 -503 1011
rect -445 1045 -345 1061
rect -445 1011 -429 1045
rect -361 1011 -345 1045
rect -445 964 -345 1011
rect -287 1045 -187 1061
rect -287 1011 -271 1045
rect -203 1011 -187 1045
rect -287 964 -187 1011
rect -129 1045 -29 1061
rect -129 1011 -113 1045
rect -45 1011 -29 1045
rect -129 964 -29 1011
rect 29 1045 129 1061
rect 29 1011 45 1045
rect 113 1011 129 1045
rect 29 964 129 1011
rect 187 1045 287 1061
rect 187 1011 203 1045
rect 271 1011 287 1045
rect 187 964 287 1011
rect 345 1045 445 1061
rect 345 1011 361 1045
rect 429 1011 445 1045
rect 345 964 445 1011
rect 503 1045 603 1061
rect 503 1011 519 1045
rect 587 1011 603 1045
rect 503 964 603 1011
rect 661 1045 761 1061
rect 661 1011 677 1045
rect 745 1011 761 1045
rect 661 964 761 1011
rect -761 -1062 -661 -1036
rect -603 -1062 -503 -1036
rect -445 -1062 -345 -1036
rect -287 -1062 -187 -1036
rect -129 -1062 -29 -1036
rect 29 -1062 129 -1036
rect 187 -1062 287 -1036
rect 345 -1062 445 -1036
rect 503 -1062 603 -1036
rect 661 -1062 761 -1036
<< polycont >>
rect -745 1011 -677 1045
rect -587 1011 -519 1045
rect -429 1011 -361 1045
rect -271 1011 -203 1045
rect -113 1011 -45 1045
rect 45 1011 113 1045
rect 203 1011 271 1045
rect 361 1011 429 1045
rect 519 1011 587 1045
rect 677 1011 745 1045
<< locali >>
rect -761 1011 -745 1045
rect -677 1011 -661 1045
rect -603 1011 -587 1045
rect -519 1011 -503 1045
rect -445 1011 -429 1045
rect -361 1011 -345 1045
rect -287 1011 -271 1045
rect -203 1011 -187 1045
rect -129 1011 -113 1045
rect -45 1011 -29 1045
rect 29 1011 45 1045
rect 113 1011 129 1045
rect 187 1011 203 1045
rect 271 1011 287 1045
rect 345 1011 361 1045
rect 429 1011 445 1045
rect 503 1011 519 1045
rect 587 1011 603 1045
rect 661 1011 677 1045
rect 745 1011 761 1045
rect -807 952 -773 968
rect -807 -1040 -773 -1024
rect -649 952 -615 968
rect -649 -1040 -615 -1024
rect -491 952 -457 968
rect -491 -1040 -457 -1024
rect -333 952 -299 968
rect -333 -1040 -299 -1024
rect -175 952 -141 968
rect -175 -1040 -141 -1024
rect -17 952 17 968
rect -17 -1040 17 -1024
rect 141 952 175 968
rect 141 -1040 175 -1024
rect 299 952 333 968
rect 299 -1040 333 -1024
rect 457 952 491 968
rect 457 -1040 491 -1024
rect 615 952 649 968
rect 615 -1040 649 -1024
rect 773 952 807 968
rect 773 -1040 807 -1024
<< viali >>
rect -745 1011 -677 1045
rect -587 1011 -519 1045
rect -429 1011 -361 1045
rect -271 1011 -203 1045
rect -113 1011 -45 1045
rect 45 1011 113 1045
rect 203 1011 271 1045
rect 361 1011 429 1045
rect 519 1011 587 1045
rect 677 1011 745 1045
rect -807 -1007 -773 -414
rect -649 342 -615 935
rect -491 -1007 -457 -414
rect -333 342 -299 935
rect -175 -1007 -141 -414
rect -17 342 17 935
rect 141 -1007 175 -414
rect 299 342 333 935
rect 457 -1007 491 -414
rect 615 342 649 935
rect 773 -1007 807 -414
<< metal1 >>
rect -757 1045 -665 1051
rect -757 1011 -745 1045
rect -677 1011 -665 1045
rect -757 1005 -665 1011
rect -599 1045 -507 1051
rect -599 1011 -587 1045
rect -519 1011 -507 1045
rect -599 1005 -507 1011
rect -441 1045 -349 1051
rect -441 1011 -429 1045
rect -361 1011 -349 1045
rect -441 1005 -349 1011
rect -283 1045 -191 1051
rect -283 1011 -271 1045
rect -203 1011 -191 1045
rect -283 1005 -191 1011
rect -125 1045 -33 1051
rect -125 1011 -113 1045
rect -45 1011 -33 1045
rect -125 1005 -33 1011
rect 33 1045 125 1051
rect 33 1011 45 1045
rect 113 1011 125 1045
rect 33 1005 125 1011
rect 191 1045 283 1051
rect 191 1011 203 1045
rect 271 1011 283 1045
rect 191 1005 283 1011
rect 349 1045 441 1051
rect 349 1011 361 1045
rect 429 1011 441 1045
rect 349 1005 441 1011
rect 507 1045 599 1051
rect 507 1011 519 1045
rect 587 1011 599 1045
rect 507 1005 599 1011
rect 665 1045 757 1051
rect 665 1011 677 1045
rect 745 1011 757 1045
rect 665 1005 757 1011
rect -655 935 -609 947
rect -655 342 -649 935
rect -615 342 -609 935
rect -655 330 -609 342
rect -339 935 -293 947
rect -339 342 -333 935
rect -299 342 -293 935
rect -339 330 -293 342
rect -23 935 23 947
rect -23 342 -17 935
rect 17 342 23 935
rect -23 330 23 342
rect 293 935 339 947
rect 293 342 299 935
rect 333 342 339 935
rect 293 330 339 342
rect 609 935 655 947
rect 609 342 615 935
rect 649 342 655 935
rect 609 330 655 342
rect -813 -414 -767 -402
rect -813 -1007 -807 -414
rect -773 -1007 -767 -414
rect -813 -1019 -767 -1007
rect -497 -414 -451 -402
rect -497 -1007 -491 -414
rect -457 -1007 -451 -414
rect -497 -1019 -451 -1007
rect -181 -414 -135 -402
rect -181 -1007 -175 -414
rect -141 -1007 -135 -414
rect -181 -1019 -135 -1007
rect 135 -414 181 -402
rect 135 -1007 141 -414
rect 175 -1007 181 -414
rect 135 -1019 181 -1007
rect 451 -414 497 -402
rect 451 -1007 457 -414
rect 491 -1007 497 -414
rect 451 -1019 497 -1007
rect 767 -414 813 -402
rect 767 -1007 773 -414
rect 807 -1007 813 -414
rect 767 -1019 813 -1007
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc -30 viadrn +30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
