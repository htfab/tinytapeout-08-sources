magic
tech sky130A
timestamp 1725574488
<< metal1 >>
rect 5900 5545 6000 5645
rect 6385 5545 6485 5645
rect 9445 5545 9545 5645
rect 9935 5545 10035 5645
rect 3265 1850 3900 1950
rect 3265 1755 3720 1760
rect 3265 1685 3655 1755
rect 3715 1685 3720 1755
rect 3265 1660 3720 1685
rect 3505 1545 3600 1550
rect 3505 1465 3510 1545
rect 3595 1465 3600 1545
rect 3505 1460 3600 1465
rect 3505 -3330 3575 1460
rect 3650 -2800 3720 1660
rect 5895 -2205 5995 -2105
rect 6385 -2205 6485 -2105
rect 9445 -2205 9545 -2105
rect 9935 -2205 10035 -2105
rect 3945 -2715 5285 -2710
rect 3945 -2770 3950 -2715
rect 4065 -2770 5285 -2715
rect 3945 -2775 5285 -2770
rect 5190 -2800 5285 -2775
rect 5585 -2800 5685 -2685
rect 3650 -2900 3800 -2800
rect 3505 -3430 3900 -3330
rect 4620 -3825 4720 -3430
rect 5190 -3825 5290 -3430
<< via1 >>
rect 3655 1685 3715 1755
rect 4550 1685 4680 1755
rect 3510 1465 3595 1545
rect 4400 1455 4495 1545
rect 3980 -1775 4040 -1690
rect 3950 -2770 4065 -2715
<< metal2 >>
rect 3650 1755 4685 1760
rect 3650 1685 3655 1755
rect 3715 1685 4550 1755
rect 4680 1685 4685 1755
rect 3650 1680 4685 1685
rect 3505 1545 3600 1550
rect 3505 1465 3510 1545
rect 3595 1530 3600 1545
rect 4395 1545 4500 1550
rect 4395 1530 4400 1545
rect 3595 1475 4400 1530
rect 3595 1465 3600 1475
rect 3505 1460 3600 1465
rect 4395 1455 4400 1475
rect 4495 1455 4500 1545
rect 4395 1450 4500 1455
rect 3975 -1690 4045 -1685
rect 3975 -1775 3980 -1690
rect 4040 -1775 4045 -1690
rect 3975 -2710 4045 -1775
rect 3945 -2715 4070 -2710
rect 3945 -2770 3950 -2715
rect 4065 -2770 4070 -2715
rect 3945 -2775 4070 -2770
use vco_bias  x1
timestamp 1725572295
transform 1 0 3540 0 -1 -3330
box 260 -530 2145 100
use vco_core  x6
timestamp 1725572295
transform 1 0 5100 0 1 2390
box -1300 -5080 7005 3740
<< labels >>
flabel metal1 3265 1850 3365 1950 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel metal1 3265 1660 3365 1760 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel metal1 4620 -3825 4720 -3725 0 FreeSans 640 0 0 0 Icont
port 2 nsew
flabel metal1 5190 -3825 5290 -3725 0 FreeSans 640 0 0 0 Vb
port 11 nsew
flabel metal1 5900 5545 6000 5645 0 FreeSans 640 0 0 0 Vp0
port 3 nsew
flabel metal1 6385 5545 6485 5645 0 FreeSans 640 0 0 0 Vn0
port 7 nsew
flabel metal1 9935 5545 10035 5645 0 FreeSans 640 0 0 0 Vp1
port 4 nsew
flabel metal1 9445 5545 9545 5645 0 FreeSans 640 0 0 0 Vn1
port 8 nsew
flabel metal1 9935 -2205 10035 -2105 0 FreeSans 640 0 0 0 Vp2
port 5 nsew
flabel metal1 9445 -2205 9545 -2105 0 FreeSans 640 0 0 0 Vn2
port 9 nsew
flabel metal1 5895 -2205 5995 -2105 0 FreeSans 640 0 0 0 Vp3
port 6 nsew
flabel metal1 6385 -2205 6485 -2105 0 FreeSans 640 0 0 0 Vn3
port 10 nsew
<< end >>
