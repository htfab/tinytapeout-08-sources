magic
tech sky130A
magscale 1 2
timestamp 1725402679
<< nwell >>
rect -1803 -498 1803 464
<< pmoslvt >>
rect -1709 -436 -1609 364
rect -1551 -436 -1451 364
rect -1393 -436 -1293 364
rect -1235 -436 -1135 364
rect -1077 -436 -977 364
rect -919 -436 -819 364
rect -761 -436 -661 364
rect -603 -436 -503 364
rect -445 -436 -345 364
rect -287 -436 -187 364
rect -129 -436 -29 364
rect 29 -436 129 364
rect 187 -436 287 364
rect 345 -436 445 364
rect 503 -436 603 364
rect 661 -436 761 364
rect 819 -436 919 364
rect 977 -436 1077 364
rect 1135 -436 1235 364
rect 1293 -436 1393 364
rect 1451 -436 1551 364
rect 1609 -436 1709 364
<< pdiff >>
rect -1767 352 -1709 364
rect -1767 -424 -1755 352
rect -1721 -424 -1709 352
rect -1767 -436 -1709 -424
rect -1609 352 -1551 364
rect -1609 -424 -1597 352
rect -1563 -424 -1551 352
rect -1609 -436 -1551 -424
rect -1451 352 -1393 364
rect -1451 -424 -1439 352
rect -1405 -424 -1393 352
rect -1451 -436 -1393 -424
rect -1293 352 -1235 364
rect -1293 -424 -1281 352
rect -1247 -424 -1235 352
rect -1293 -436 -1235 -424
rect -1135 352 -1077 364
rect -1135 -424 -1123 352
rect -1089 -424 -1077 352
rect -1135 -436 -1077 -424
rect -977 352 -919 364
rect -977 -424 -965 352
rect -931 -424 -919 352
rect -977 -436 -919 -424
rect -819 352 -761 364
rect -819 -424 -807 352
rect -773 -424 -761 352
rect -819 -436 -761 -424
rect -661 352 -603 364
rect -661 -424 -649 352
rect -615 -424 -603 352
rect -661 -436 -603 -424
rect -503 352 -445 364
rect -503 -424 -491 352
rect -457 -424 -445 352
rect -503 -436 -445 -424
rect -345 352 -287 364
rect -345 -424 -333 352
rect -299 -424 -287 352
rect -345 -436 -287 -424
rect -187 352 -129 364
rect -187 -424 -175 352
rect -141 -424 -129 352
rect -187 -436 -129 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 129 352 187 364
rect 129 -424 141 352
rect 175 -424 187 352
rect 129 -436 187 -424
rect 287 352 345 364
rect 287 -424 299 352
rect 333 -424 345 352
rect 287 -436 345 -424
rect 445 352 503 364
rect 445 -424 457 352
rect 491 -424 503 352
rect 445 -436 503 -424
rect 603 352 661 364
rect 603 -424 615 352
rect 649 -424 661 352
rect 603 -436 661 -424
rect 761 352 819 364
rect 761 -424 773 352
rect 807 -424 819 352
rect 761 -436 819 -424
rect 919 352 977 364
rect 919 -424 931 352
rect 965 -424 977 352
rect 919 -436 977 -424
rect 1077 352 1135 364
rect 1077 -424 1089 352
rect 1123 -424 1135 352
rect 1077 -436 1135 -424
rect 1235 352 1293 364
rect 1235 -424 1247 352
rect 1281 -424 1293 352
rect 1235 -436 1293 -424
rect 1393 352 1451 364
rect 1393 -424 1405 352
rect 1439 -424 1451 352
rect 1393 -436 1451 -424
rect 1551 352 1609 364
rect 1551 -424 1563 352
rect 1597 -424 1609 352
rect 1551 -436 1609 -424
rect 1709 352 1767 364
rect 1709 -424 1721 352
rect 1755 -424 1767 352
rect 1709 -436 1767 -424
<< pdiffc >>
rect -1755 -424 -1721 352
rect -1597 -424 -1563 352
rect -1439 -424 -1405 352
rect -1281 -424 -1247 352
rect -1123 -424 -1089 352
rect -965 -424 -931 352
rect -807 -424 -773 352
rect -649 -424 -615 352
rect -491 -424 -457 352
rect -333 -424 -299 352
rect -175 -424 -141 352
rect -17 -424 17 352
rect 141 -424 175 352
rect 299 -424 333 352
rect 457 -424 491 352
rect 615 -424 649 352
rect 773 -424 807 352
rect 931 -424 965 352
rect 1089 -424 1123 352
rect 1247 -424 1281 352
rect 1405 -424 1439 352
rect 1563 -424 1597 352
rect 1721 -424 1755 352
<< poly >>
rect -1709 445 -1609 461
rect -1709 411 -1693 445
rect -1625 411 -1609 445
rect -1709 364 -1609 411
rect -1551 445 -1451 461
rect -1551 411 -1535 445
rect -1467 411 -1451 445
rect -1551 364 -1451 411
rect -1393 445 -1293 461
rect -1393 411 -1377 445
rect -1309 411 -1293 445
rect -1393 364 -1293 411
rect -1235 445 -1135 461
rect -1235 411 -1219 445
rect -1151 411 -1135 445
rect -1235 364 -1135 411
rect -1077 445 -977 461
rect -1077 411 -1061 445
rect -993 411 -977 445
rect -1077 364 -977 411
rect -919 445 -819 461
rect -919 411 -903 445
rect -835 411 -819 445
rect -919 364 -819 411
rect -761 445 -661 461
rect -761 411 -745 445
rect -677 411 -661 445
rect -761 364 -661 411
rect -603 445 -503 461
rect -603 411 -587 445
rect -519 411 -503 445
rect -603 364 -503 411
rect -445 445 -345 461
rect -445 411 -429 445
rect -361 411 -345 445
rect -445 364 -345 411
rect -287 445 -187 461
rect -287 411 -271 445
rect -203 411 -187 445
rect -287 364 -187 411
rect -129 445 -29 461
rect -129 411 -113 445
rect -45 411 -29 445
rect -129 364 -29 411
rect 29 445 129 461
rect 29 411 45 445
rect 113 411 129 445
rect 29 364 129 411
rect 187 445 287 461
rect 187 411 203 445
rect 271 411 287 445
rect 187 364 287 411
rect 345 445 445 461
rect 345 411 361 445
rect 429 411 445 445
rect 345 364 445 411
rect 503 445 603 461
rect 503 411 519 445
rect 587 411 603 445
rect 503 364 603 411
rect 661 445 761 461
rect 661 411 677 445
rect 745 411 761 445
rect 661 364 761 411
rect 819 445 919 461
rect 819 411 835 445
rect 903 411 919 445
rect 819 364 919 411
rect 977 445 1077 461
rect 977 411 993 445
rect 1061 411 1077 445
rect 977 364 1077 411
rect 1135 445 1235 461
rect 1135 411 1151 445
rect 1219 411 1235 445
rect 1135 364 1235 411
rect 1293 445 1393 461
rect 1293 411 1309 445
rect 1377 411 1393 445
rect 1293 364 1393 411
rect 1451 445 1551 461
rect 1451 411 1467 445
rect 1535 411 1551 445
rect 1451 364 1551 411
rect 1609 445 1709 461
rect 1609 411 1625 445
rect 1693 411 1709 445
rect 1609 364 1709 411
rect -1709 -462 -1609 -436
rect -1551 -462 -1451 -436
rect -1393 -462 -1293 -436
rect -1235 -462 -1135 -436
rect -1077 -462 -977 -436
rect -919 -462 -819 -436
rect -761 -462 -661 -436
rect -603 -462 -503 -436
rect -445 -462 -345 -436
rect -287 -462 -187 -436
rect -129 -462 -29 -436
rect 29 -462 129 -436
rect 187 -462 287 -436
rect 345 -462 445 -436
rect 503 -462 603 -436
rect 661 -462 761 -436
rect 819 -462 919 -436
rect 977 -462 1077 -436
rect 1135 -462 1235 -436
rect 1293 -462 1393 -436
rect 1451 -462 1551 -436
rect 1609 -462 1709 -436
<< polycont >>
rect -1693 411 -1625 445
rect -1535 411 -1467 445
rect -1377 411 -1309 445
rect -1219 411 -1151 445
rect -1061 411 -993 445
rect -903 411 -835 445
rect -745 411 -677 445
rect -587 411 -519 445
rect -429 411 -361 445
rect -271 411 -203 445
rect -113 411 -45 445
rect 45 411 113 445
rect 203 411 271 445
rect 361 411 429 445
rect 519 411 587 445
rect 677 411 745 445
rect 835 411 903 445
rect 993 411 1061 445
rect 1151 411 1219 445
rect 1309 411 1377 445
rect 1467 411 1535 445
rect 1625 411 1693 445
<< locali >>
rect -1709 411 -1693 445
rect -1625 411 -1609 445
rect -1551 411 -1535 445
rect -1467 411 -1451 445
rect -1393 411 -1377 445
rect -1309 411 -1293 445
rect -1235 411 -1219 445
rect -1151 411 -1135 445
rect -1077 411 -1061 445
rect -993 411 -977 445
rect -919 411 -903 445
rect -835 411 -819 445
rect -761 411 -745 445
rect -677 411 -661 445
rect -603 411 -587 445
rect -519 411 -503 445
rect -445 411 -429 445
rect -361 411 -345 445
rect -287 411 -271 445
rect -203 411 -187 445
rect -129 411 -113 445
rect -45 411 -29 445
rect 29 411 45 445
rect 113 411 129 445
rect 187 411 203 445
rect 271 411 287 445
rect 345 411 361 445
rect 429 411 445 445
rect 503 411 519 445
rect 587 411 603 445
rect 661 411 677 445
rect 745 411 761 445
rect 819 411 835 445
rect 903 411 919 445
rect 977 411 993 445
rect 1061 411 1077 445
rect 1135 411 1151 445
rect 1219 411 1235 445
rect 1293 411 1309 445
rect 1377 411 1393 445
rect 1451 411 1467 445
rect 1535 411 1551 445
rect 1609 411 1625 445
rect 1693 411 1709 445
rect -1755 352 -1721 368
rect -1755 -440 -1721 -424
rect -1597 352 -1563 368
rect -1597 -440 -1563 -424
rect -1439 352 -1405 368
rect -1439 -440 -1405 -424
rect -1281 352 -1247 368
rect -1281 -440 -1247 -424
rect -1123 352 -1089 368
rect -1123 -440 -1089 -424
rect -965 352 -931 368
rect -965 -440 -931 -424
rect -807 352 -773 368
rect -807 -440 -773 -424
rect -649 352 -615 368
rect -649 -440 -615 -424
rect -491 352 -457 368
rect -491 -440 -457 -424
rect -333 352 -299 368
rect -333 -440 -299 -424
rect -175 352 -141 368
rect -175 -440 -141 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 141 352 175 368
rect 141 -440 175 -424
rect 299 352 333 368
rect 299 -440 333 -424
rect 457 352 491 368
rect 457 -440 491 -424
rect 615 352 649 368
rect 615 -440 649 -424
rect 773 352 807 368
rect 773 -440 807 -424
rect 931 352 965 368
rect 931 -440 965 -424
rect 1089 352 1123 368
rect 1089 -440 1123 -424
rect 1247 352 1281 368
rect 1247 -440 1281 -424
rect 1405 352 1439 368
rect 1405 -440 1439 -424
rect 1563 352 1597 368
rect 1563 -440 1597 -424
rect 1721 352 1755 368
rect 1721 -440 1755 -424
<< viali >>
rect -1693 411 -1625 445
rect -1535 411 -1467 445
rect -1377 411 -1309 445
rect -1219 411 -1151 445
rect -1061 411 -993 445
rect -903 411 -835 445
rect -745 411 -677 445
rect -587 411 -519 445
rect -429 411 -361 445
rect -271 411 -203 445
rect -113 411 -45 445
rect 45 411 113 445
rect 203 411 271 445
rect 361 411 429 445
rect 519 411 587 445
rect 677 411 745 445
rect 835 411 903 445
rect 993 411 1061 445
rect 1151 411 1219 445
rect 1309 411 1377 445
rect 1467 411 1535 445
rect 1625 411 1693 445
rect -1755 -407 -1721 -174
rect -1597 102 -1563 335
rect -1439 -407 -1405 -174
rect -1281 102 -1247 335
rect -1123 -407 -1089 -174
rect -965 102 -931 335
rect -807 -407 -773 -174
rect -649 102 -615 335
rect -491 -407 -457 -174
rect -333 102 -299 335
rect -175 -407 -141 -174
rect -17 102 17 335
rect 141 -407 175 -174
rect 299 102 333 335
rect 457 -407 491 -174
rect 615 102 649 335
rect 773 -407 807 -174
rect 931 102 965 335
rect 1089 -407 1123 -174
rect 1247 102 1281 335
rect 1405 -407 1439 -174
rect 1563 102 1597 335
rect 1721 -407 1755 -174
<< metal1 >>
rect -1705 445 -1613 451
rect -1705 411 -1693 445
rect -1625 411 -1613 445
rect -1705 405 -1613 411
rect -1547 445 -1455 451
rect -1547 411 -1535 445
rect -1467 411 -1455 445
rect -1547 405 -1455 411
rect -1389 445 -1297 451
rect -1389 411 -1377 445
rect -1309 411 -1297 445
rect -1389 405 -1297 411
rect -1231 445 -1139 451
rect -1231 411 -1219 445
rect -1151 411 -1139 445
rect -1231 405 -1139 411
rect -1073 445 -981 451
rect -1073 411 -1061 445
rect -993 411 -981 445
rect -1073 405 -981 411
rect -915 445 -823 451
rect -915 411 -903 445
rect -835 411 -823 445
rect -915 405 -823 411
rect -757 445 -665 451
rect -757 411 -745 445
rect -677 411 -665 445
rect -757 405 -665 411
rect -599 445 -507 451
rect -599 411 -587 445
rect -519 411 -507 445
rect -599 405 -507 411
rect -441 445 -349 451
rect -441 411 -429 445
rect -361 411 -349 445
rect -441 405 -349 411
rect -283 445 -191 451
rect -283 411 -271 445
rect -203 411 -191 445
rect -283 405 -191 411
rect -125 445 -33 451
rect -125 411 -113 445
rect -45 411 -33 445
rect -125 405 -33 411
rect 33 445 125 451
rect 33 411 45 445
rect 113 411 125 445
rect 33 405 125 411
rect 191 445 283 451
rect 191 411 203 445
rect 271 411 283 445
rect 191 405 283 411
rect 349 445 441 451
rect 349 411 361 445
rect 429 411 441 445
rect 349 405 441 411
rect 507 445 599 451
rect 507 411 519 445
rect 587 411 599 445
rect 507 405 599 411
rect 665 445 757 451
rect 665 411 677 445
rect 745 411 757 445
rect 665 405 757 411
rect 823 445 915 451
rect 823 411 835 445
rect 903 411 915 445
rect 823 405 915 411
rect 981 445 1073 451
rect 981 411 993 445
rect 1061 411 1073 445
rect 981 405 1073 411
rect 1139 445 1231 451
rect 1139 411 1151 445
rect 1219 411 1231 445
rect 1139 405 1231 411
rect 1297 445 1389 451
rect 1297 411 1309 445
rect 1377 411 1389 445
rect 1297 405 1389 411
rect 1455 445 1547 451
rect 1455 411 1467 445
rect 1535 411 1547 445
rect 1455 405 1547 411
rect 1613 445 1705 451
rect 1613 411 1625 445
rect 1693 411 1705 445
rect 1613 405 1705 411
rect -1603 335 -1557 347
rect -1603 102 -1597 335
rect -1563 102 -1557 335
rect -1603 90 -1557 102
rect -1287 335 -1241 347
rect -1287 102 -1281 335
rect -1247 102 -1241 335
rect -1287 90 -1241 102
rect -971 335 -925 347
rect -971 102 -965 335
rect -931 102 -925 335
rect -971 90 -925 102
rect -655 335 -609 347
rect -655 102 -649 335
rect -615 102 -609 335
rect -655 90 -609 102
rect -339 335 -293 347
rect -339 102 -333 335
rect -299 102 -293 335
rect -339 90 -293 102
rect -23 335 23 347
rect -23 102 -17 335
rect 17 102 23 335
rect -23 90 23 102
rect 293 335 339 347
rect 293 102 299 335
rect 333 102 339 335
rect 293 90 339 102
rect 609 335 655 347
rect 609 102 615 335
rect 649 102 655 335
rect 609 90 655 102
rect 925 335 971 347
rect 925 102 931 335
rect 965 102 971 335
rect 925 90 971 102
rect 1241 335 1287 347
rect 1241 102 1247 335
rect 1281 102 1287 335
rect 1241 90 1287 102
rect 1557 335 1603 347
rect 1557 102 1563 335
rect 1597 102 1603 335
rect 1557 90 1603 102
rect -1761 -174 -1715 -162
rect -1761 -407 -1755 -174
rect -1721 -407 -1715 -174
rect -1761 -419 -1715 -407
rect -1445 -174 -1399 -162
rect -1445 -407 -1439 -174
rect -1405 -407 -1399 -174
rect -1445 -419 -1399 -407
rect -1129 -174 -1083 -162
rect -1129 -407 -1123 -174
rect -1089 -407 -1083 -174
rect -1129 -419 -1083 -407
rect -813 -174 -767 -162
rect -813 -407 -807 -174
rect -773 -407 -767 -174
rect -813 -419 -767 -407
rect -497 -174 -451 -162
rect -497 -407 -491 -174
rect -457 -407 -451 -174
rect -497 -419 -451 -407
rect -181 -174 -135 -162
rect -181 -407 -175 -174
rect -141 -407 -135 -174
rect -181 -419 -135 -407
rect 135 -174 181 -162
rect 135 -407 141 -174
rect 175 -407 181 -174
rect 135 -419 181 -407
rect 451 -174 497 -162
rect 451 -407 457 -174
rect 491 -407 497 -174
rect 451 -419 497 -407
rect 767 -174 813 -162
rect 767 -407 773 -174
rect 807 -407 813 -174
rect 767 -419 813 -407
rect 1083 -174 1129 -162
rect 1083 -407 1089 -174
rect 1123 -407 1129 -174
rect 1083 -419 1129 -407
rect 1399 -174 1445 -162
rect 1399 -407 1405 -174
rect 1439 -407 1445 -174
rect 1399 -419 1445 -407
rect 1715 -174 1761 -162
rect 1715 -407 1721 -174
rect 1755 -407 1761 -174
rect 1715 -419 1761 -407
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 0.5 m 1 nf 22 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc -30 viadrn +30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
