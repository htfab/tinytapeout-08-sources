magic
tech sky130A
magscale 1 2
timestamp 1724347750
<< viali >>
rect 1758 1344 2206 1416
rect 1680 -866 2304 -822
<< metal1 >>
rect -643 2287 2201 2729
rect 621 2027 1063 2287
rect 1759 2180 2201 2287
rect 615 1585 621 2027
rect 1063 1585 1069 2027
rect 120 1306 1152 1436
rect 1736 1416 2226 2180
rect 1736 1344 1758 1416
rect 2206 1344 2226 1416
rect 1736 1336 2226 1344
rect 120 1244 2494 1306
rect 120 1236 1152 1244
rect 120 586 320 1236
rect 622 1136 1062 1142
rect 1400 1136 1476 1194
rect 1062 696 1476 1136
rect 622 690 1062 696
rect 1400 612 1476 696
rect 2504 1142 2570 1178
rect 2504 994 2732 1142
rect 2504 766 3092 994
rect 2504 634 2732 766
rect 120 578 1252 586
rect 120 509 2568 578
rect 115 386 2568 509
rect 115 366 309 386
rect 1230 378 2568 386
rect -476 174 309 366
rect -476 166 -284 174
rect 115 136 309 174
rect 2864 348 3092 766
rect 2864 148 3424 348
rect 115 -58 2580 136
rect 115 -715 309 -58
rect 1414 -128 1470 -96
rect 634 -188 1006 -182
rect 1098 -188 1470 -128
rect 628 -560 634 -188
rect 1006 -560 1470 -188
rect 634 -566 1006 -560
rect 1098 -642 1470 -560
rect 1414 -686 1470 -642
rect 2498 -304 2576 -106
rect 2864 -304 3092 148
rect 2498 -532 3092 -304
rect 2498 -684 2576 -532
rect 115 -716 1175 -715
rect 115 -718 1286 -716
rect 115 -780 2514 -718
rect 115 -792 1286 -780
rect 115 -909 1200 -792
rect 1662 -822 2324 -810
rect 1662 -866 1680 -822
rect 2304 -866 2324 -822
rect 1662 -876 2324 -866
rect 1124 -910 1200 -909
rect 1666 -1066 2312 -876
rect 628 -1448 634 -1076
rect 1006 -1448 1012 -1076
rect 634 -1538 1006 -1448
rect 1798 -1538 2170 -1066
rect 634 -1548 2170 -1538
rect -604 -1910 2170 -1548
rect -604 -1920 1006 -1910
<< via1 >>
rect 621 1585 1063 2027
rect 622 696 1062 1136
rect 634 -560 1006 -188
rect 634 -1448 1006 -1076
<< metal2 >>
rect 621 2027 1063 2033
rect 621 1136 1063 1585
rect 616 696 622 1136
rect 1062 696 1068 1136
rect 621 695 1063 696
rect 628 -560 634 -188
rect 1006 -560 1012 -188
rect 634 -1076 1006 -560
rect 634 -1454 1006 -1448
use sky130_fd_pr__nfet_01v8_Q3BYGR  XM1
timestamp 1724342599
transform 1 0 1986 0 1 -388
box -696 -510 696 510
use sky130_fd_pr__pfet_01v8_SKN7VM  XM2
timestamp 1724342599
transform 1 0 1986 0 1 907
box -696 -519 696 519
<< labels >>
flabel metal1 3224 148 3424 348 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel space -476 166 -276 366 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 -540 2390 -340 2590 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -534 -1846 -334 -1646 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
