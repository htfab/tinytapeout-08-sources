magic
tech sky130A
magscale 1 2
timestamp 1725256412
<< locali >>
rect 2868 631 3056 656
rect 2868 597 2873 631
rect 2907 597 2945 631
rect 2979 597 3017 631
rect 3051 597 3056 631
rect 2868 572 3056 597
rect 3642 623 3830 648
rect 3642 589 3647 623
rect 3681 589 3719 623
rect 3753 589 3791 623
rect 3825 589 3830 623
rect 3642 564 3830 589
rect 4408 629 4596 654
rect 4408 595 4413 629
rect 4447 595 4485 629
rect 4519 595 4557 629
rect 4591 595 4596 629
rect 4408 570 4596 595
rect 1452 -3739 1802 -3736
rect 1452 -3845 1466 -3739
rect 1788 -3845 1802 -3739
rect 1452 -3848 1802 -3845
rect -792 -4620 746 -4604
rect -792 -4726 -760 -4620
rect 714 -4726 746 -4620
rect -792 -4742 746 -4726
rect 4124 -4690 4362 -4660
rect 4124 -5156 4154 -4690
rect 4332 -5156 4362 -4690
rect 4124 -5186 4362 -5156
rect 454 -5233 784 -5206
rect 454 -5267 458 -5233
rect 492 -5267 530 -5233
rect 564 -5267 602 -5233
rect 636 -5267 674 -5233
rect 708 -5267 746 -5233
rect 780 -5267 784 -5233
rect 454 -5294 784 -5267
rect 1568 -5264 1806 -5232
rect 1568 -5298 1598 -5264
rect 1632 -5298 1670 -5264
rect 1704 -5298 1742 -5264
rect 1776 -5298 1806 -5264
rect 1568 -5330 1806 -5298
rect 3008 -5262 3292 -5238
rect 3008 -5296 3025 -5262
rect 3059 -5296 3097 -5262
rect 3131 -5296 3169 -5262
rect 3203 -5296 3241 -5262
rect 3275 -5296 3292 -5262
rect 3008 -5320 3292 -5296
rect 4112 -5259 4288 -5246
rect 4112 -5365 4147 -5259
rect 4253 -5365 4288 -5259
rect 4112 -5378 4288 -5365
<< viali >>
rect 2873 597 2907 631
rect 2945 597 2979 631
rect 3017 597 3051 631
rect 3647 589 3681 623
rect 3719 589 3753 623
rect 3791 589 3825 623
rect 4413 595 4447 629
rect 4485 595 4519 629
rect 4557 595 4591 629
rect 1466 -3845 1788 -3739
rect -760 -4726 714 -4620
rect 4154 -5156 4332 -4690
rect 458 -5267 492 -5233
rect 530 -5267 564 -5233
rect 602 -5267 636 -5233
rect 674 -5267 708 -5233
rect 746 -5267 780 -5233
rect 1598 -5298 1632 -5264
rect 1670 -5298 1704 -5264
rect 1742 -5298 1776 -5264
rect 3025 -5296 3059 -5262
rect 3097 -5296 3131 -5262
rect 3169 -5296 3203 -5262
rect 3241 -5296 3275 -5262
rect 4147 -5365 4253 -5259
<< metal1 >>
rect -1102 660 4596 1024
rect -1102 640 4608 660
rect -1102 588 2872 640
rect 2924 588 2936 640
rect 2988 588 3000 640
rect 3052 638 4608 640
rect 3052 632 4412 638
rect 3052 588 3646 632
rect -1102 580 3646 588
rect 3698 580 3710 632
rect 3762 580 3774 632
rect 3826 586 4412 632
rect 4464 586 4476 638
rect 4528 586 4540 638
rect 4592 586 4608 638
rect 3826 580 4608 586
rect -1102 564 4608 580
rect -1102 560 4596 564
rect -880 72 -702 560
rect 3630 558 3842 560
rect 2762 462 4024 530
rect 4132 512 4212 524
rect 4132 464 4706 512
rect 2796 282 2898 462
rect 3050 288 3124 462
rect 2662 199 2770 214
rect 2662 147 2690 199
rect 2742 147 2770 199
rect 2662 135 2770 147
rect 2662 83 2690 135
rect 2742 83 2770 135
rect -842 54 -746 72
rect 2662 68 2770 83
rect 2904 201 3012 216
rect 2904 149 2932 201
rect 2984 149 3012 201
rect 2904 137 3012 149
rect 2904 85 2932 137
rect 2984 85 3012 137
rect 2904 70 3012 85
rect 3140 195 3248 210
rect 3140 143 3168 195
rect 3220 143 3248 195
rect 3140 131 3248 143
rect 3140 79 3168 131
rect 3220 79 3248 131
rect 3140 64 3248 79
rect -380 -156 4 -20
rect 408 -130 800 -22
rect 906 -506 986 -498
rect 1822 -506 2318 -504
rect 906 -570 1482 -506
rect 1822 -562 2322 -506
rect -1268 -1790 -1148 -1774
rect -1268 -1800 -1234 -1790
rect -1366 -1842 -1234 -1800
rect -1182 -1800 -1148 -1790
rect -1182 -1842 -1106 -1800
rect -1366 -1854 -1106 -1842
rect -1366 -1906 -1234 -1854
rect -1182 -1906 -1106 -1854
rect -1366 -1918 -1106 -1906
rect -1366 -1970 -1234 -1918
rect -1182 -1970 -1106 -1918
rect -1366 -1982 -1106 -1970
rect -1366 -2000 -1234 -1982
rect -1268 -2034 -1234 -2000
rect -1182 -2000 -1106 -1982
rect -1182 -2034 -1148 -2000
rect -1268 -2050 -1148 -2034
rect -1418 -2649 -1064 -2558
rect 906 -2646 986 -570
rect 1330 -901 1434 -876
rect 1330 -953 1356 -901
rect 1408 -953 1434 -901
rect 1330 -965 1434 -953
rect 1330 -1017 1356 -965
rect 1408 -1017 1434 -965
rect 1330 -1029 1434 -1017
rect 1330 -1081 1356 -1029
rect 1408 -1081 1434 -1029
rect 1330 -1093 1434 -1081
rect 1330 -1145 1356 -1093
rect 1408 -1145 1434 -1093
rect 1330 -1170 1434 -1145
rect 2248 -1694 2322 -562
rect 2800 -903 2904 -878
rect 2800 -955 2826 -903
rect 2878 -955 2904 -903
rect 2800 -967 2904 -955
rect 2800 -1019 2826 -967
rect 2878 -1019 2904 -967
rect 2800 -1031 2904 -1019
rect 2800 -1083 2826 -1031
rect 2878 -1083 2904 -1031
rect 2800 -1095 2904 -1083
rect 2800 -1147 2826 -1095
rect 2878 -1147 2904 -1095
rect 2800 -1172 2904 -1147
rect 3034 -903 3138 -878
rect 3034 -955 3060 -903
rect 3112 -955 3138 -903
rect 3034 -967 3138 -955
rect 3034 -1019 3060 -967
rect 3112 -1019 3138 -967
rect 3034 -1031 3138 -1019
rect 3034 -1083 3060 -1031
rect 3112 -1083 3138 -1031
rect 3034 -1095 3138 -1083
rect 3034 -1147 3060 -1095
rect 3112 -1147 3138 -1095
rect 3034 -1172 3138 -1147
rect 2220 -1708 2340 -1694
rect 2220 -1760 2254 -1708
rect 2306 -1760 2340 -1708
rect 2220 -1772 2340 -1760
rect 2220 -1824 2254 -1772
rect 2306 -1824 2340 -1772
rect 2220 -1836 2340 -1824
rect 2220 -1888 2254 -1836
rect 2306 -1888 2340 -1836
rect 2220 -1900 2340 -1888
rect 2220 -1952 2254 -1900
rect 2306 -1952 2340 -1900
rect 2220 -1966 2340 -1952
rect 1892 -2228 1992 -2198
rect 1892 -2280 1916 -2228
rect 1968 -2280 1992 -2228
rect 1892 -2292 1992 -2280
rect 1892 -2344 1916 -2292
rect 1968 -2344 1992 -2292
rect 1892 -2356 1992 -2344
rect 1892 -2408 1916 -2356
rect 1968 -2408 1992 -2356
rect 1892 -2438 1992 -2408
rect -1418 -2829 -1306 -2649
rect -1190 -2829 -1064 -2649
rect -1418 -2912 -1064 -2829
rect 872 -2675 1012 -2646
rect 872 -2855 884 -2675
rect 1000 -2855 1012 -2675
rect 872 -2884 1012 -2855
rect 906 -3630 986 -2884
rect 1200 -3364 1308 -3336
rect 1200 -3416 1228 -3364
rect 1280 -3416 1308 -3364
rect 1200 -3428 1308 -3416
rect 1200 -3480 1228 -3428
rect 1280 -3480 1308 -3428
rect 1200 -3508 1308 -3480
rect 1434 -3372 1542 -3344
rect 1434 -3424 1462 -3372
rect 1514 -3424 1542 -3372
rect 1434 -3436 1542 -3424
rect 1434 -3488 1462 -3436
rect 1514 -3488 1542 -3436
rect 1434 -3516 1542 -3488
rect 1774 -3365 1866 -3340
rect 1774 -3417 1794 -3365
rect 1846 -3417 1866 -3365
rect 1774 -3429 1866 -3417
rect 1774 -3481 1794 -3429
rect 1846 -3481 1866 -3429
rect 1774 -3506 1866 -3481
rect 2016 -3367 2108 -3342
rect 2016 -3419 2036 -3367
rect 2088 -3419 2108 -3367
rect 2016 -3431 2108 -3419
rect 2016 -3483 2036 -3431
rect 2088 -3483 2108 -3431
rect 2016 -3508 2108 -3483
rect 2248 -3630 2322 -1966
rect 2810 -2614 2884 -2478
rect 3044 -2614 3118 -2462
rect 3310 -2614 3408 462
rect 3468 191 3576 206
rect 3468 139 3496 191
rect 3548 139 3576 191
rect 3468 127 3576 139
rect 3468 75 3496 127
rect 3548 75 3576 127
rect 3468 60 3576 75
rect 3708 181 3816 196
rect 3708 129 3736 181
rect 3788 129 3816 181
rect 3708 117 3816 129
rect 3708 65 3736 117
rect 3788 65 3816 117
rect 3708 50 3816 65
rect 3946 175 4054 190
rect 3946 123 3974 175
rect 4026 123 4054 175
rect 3946 111 4054 123
rect 3946 59 3974 111
rect 4026 59 4054 111
rect 3946 44 4054 59
rect 3596 -2226 3696 -2196
rect 4132 -2198 4212 464
rect 4268 175 4376 190
rect 4268 123 4296 175
rect 4348 123 4376 175
rect 4268 111 4376 123
rect 4268 59 4296 111
rect 4348 59 4376 111
rect 4268 44 4376 59
rect 4482 181 4576 194
rect 4482 129 4503 181
rect 4555 129 4576 181
rect 4482 117 4576 129
rect 4482 65 4503 117
rect 4555 65 4576 117
rect 4482 52 4576 65
rect 4678 185 4772 198
rect 4678 133 4699 185
rect 4751 133 4772 185
rect 4678 121 4772 133
rect 4678 69 4699 121
rect 4751 69 4772 121
rect 4678 56 4772 69
rect 3596 -2278 3620 -2226
rect 3672 -2278 3696 -2226
rect 3596 -2290 3696 -2278
rect 3596 -2342 3620 -2290
rect 3672 -2342 3696 -2290
rect 3596 -2354 3696 -2342
rect 3596 -2406 3620 -2354
rect 3672 -2406 3696 -2354
rect 3596 -2436 3696 -2406
rect 3830 -2232 3930 -2202
rect 3830 -2284 3854 -2232
rect 3906 -2284 3930 -2232
rect 3830 -2296 3930 -2284
rect 3830 -2348 3854 -2296
rect 3906 -2348 3930 -2296
rect 3830 -2360 3930 -2348
rect 3830 -2412 3854 -2360
rect 3906 -2412 3930 -2360
rect 3830 -2442 3930 -2412
rect 4120 -2227 4220 -2198
rect 4120 -2279 4144 -2227
rect 4196 -2279 4220 -2227
rect 4120 -2291 4220 -2279
rect 4120 -2343 4144 -2291
rect 4196 -2343 4220 -2291
rect 4120 -2355 4220 -2343
rect 4120 -2407 4144 -2355
rect 4196 -2407 4220 -2355
rect 4120 -2436 4220 -2407
rect 2740 -2674 4012 -2614
rect 2420 -3006 2520 -2990
rect 2420 -3072 3712 -3006
rect 906 -3690 1476 -3630
rect 906 -3700 986 -3690
rect 1836 -3706 2332 -3630
rect 1440 -3739 1814 -3730
rect 1440 -3845 1466 -3739
rect 1788 -3845 1814 -3739
rect 1440 -3854 1814 -3845
rect 1012 -4016 1064 -3996
rect 2420 -4008 2520 -3072
rect 2882 -3204 3014 -3188
rect 2882 -3256 2922 -3204
rect 2974 -3256 3014 -3204
rect 2882 -3268 3014 -3256
rect 2882 -3320 2922 -3268
rect 2974 -3320 3014 -3268
rect 2882 -3336 3014 -3320
rect 3398 -3216 3530 -3200
rect 3398 -3268 3438 -3216
rect 3490 -3268 3530 -3216
rect 3398 -3280 3530 -3268
rect 3398 -3332 3438 -3280
rect 3490 -3332 3530 -3280
rect 3398 -3348 3530 -3332
rect 4132 -3418 4212 -2436
rect 13048 -2718 14714 -2692
rect 4388 -3203 4474 -3186
rect 4388 -3255 4405 -3203
rect 4457 -3255 4474 -3203
rect 4388 -3267 4474 -3255
rect 4388 -3319 4405 -3267
rect 4457 -3319 4474 -3267
rect 4388 -3336 4474 -3319
rect 4584 -3201 4670 -3184
rect 4584 -3253 4601 -3201
rect 4653 -3253 4670 -3201
rect 4584 -3265 4670 -3253
rect 4584 -3317 4601 -3265
rect 4653 -3317 4670 -3265
rect 4584 -3334 4670 -3317
rect 4120 -3466 4662 -3418
rect 4132 -3470 4340 -3466
rect 2218 -4016 2520 -4008
rect 1012 -4064 2520 -4016
rect 1012 -4066 2240 -4064
rect 1012 -4248 1064 -4066
rect -790 -4412 -406 -4276
rect 22 -4418 406 -4282
rect 802 -4378 1064 -4248
rect 1420 -4161 1544 -4144
rect 1420 -4213 1456 -4161
rect 1508 -4213 1544 -4161
rect 1420 -4225 1544 -4213
rect 1420 -4277 1456 -4225
rect 1508 -4277 1544 -4225
rect 1420 -4294 1544 -4277
rect 1938 -4161 2062 -4144
rect 1938 -4213 1974 -4161
rect 2026 -4213 2062 -4161
rect 1938 -4225 2062 -4213
rect 1938 -4277 1974 -4225
rect 2026 -4277 2062 -4225
rect 1938 -4294 2062 -4277
rect -804 -4620 758 -4598
rect -804 -4726 -760 -4620
rect 714 -4726 758 -4620
rect -804 -4748 758 -4726
rect 1012 -4780 1064 -4378
rect 1012 -4782 1066 -4780
rect 388 -4806 586 -4782
rect 650 -4806 1066 -4782
rect 388 -4830 1066 -4806
rect 388 -4840 830 -4830
rect 832 -4838 1066 -4830
rect 286 -4903 398 -4902
rect 286 -4955 316 -4903
rect 368 -4955 398 -4903
rect 576 -4936 666 -4840
rect 818 -4927 930 -4918
rect 286 -4967 398 -4955
rect 286 -5019 316 -4967
rect 368 -5019 398 -4967
rect 286 -5031 398 -5019
rect 286 -5083 316 -5031
rect 368 -5083 398 -5031
rect 818 -4979 848 -4927
rect 900 -4979 930 -4927
rect 818 -4991 930 -4979
rect 818 -5043 848 -4991
rect 900 -5043 930 -4991
rect 818 -5052 930 -5043
rect 286 -5084 398 -5083
rect 1012 -5112 1066 -4838
rect 1170 -4947 1294 -4930
rect 1170 -4999 1206 -4947
rect 1258 -4999 1294 -4947
rect 1170 -5011 1294 -4999
rect 1170 -5063 1206 -5011
rect 1258 -5063 1294 -5011
rect 1170 -5080 1294 -5063
rect 1680 -4957 1804 -4940
rect 1680 -5009 1716 -4957
rect 1768 -5009 1804 -4957
rect 1680 -5021 1804 -5009
rect 1680 -5073 1716 -5021
rect 1768 -5073 1804 -5021
rect 1680 -5090 1804 -5073
rect 2192 -4961 2316 -4944
rect 2192 -5013 2228 -4961
rect 2280 -5013 2316 -4961
rect 2192 -5025 2316 -5013
rect 2192 -5077 2228 -5025
rect 2280 -5077 2316 -5025
rect 2192 -5094 2316 -5077
rect 388 -5130 1066 -5112
rect 388 -5132 2238 -5130
rect 2420 -5132 2520 -4064
rect 4138 -4234 4340 -3470
rect 13048 -3602 13087 -2718
rect 14675 -3602 14714 -2718
rect 13048 -3628 14714 -3602
rect 4118 -4660 4368 -4648
rect 4114 -4673 4372 -4660
rect 2622 -4913 2756 -4894
rect 2622 -4965 2663 -4913
rect 2715 -4965 2756 -4913
rect 2622 -4977 2756 -4965
rect 2622 -5029 2663 -4977
rect 2715 -5029 2756 -4977
rect 2622 -5048 2756 -5029
rect 3140 -4915 3274 -4896
rect 3140 -4967 3181 -4915
rect 3233 -4967 3274 -4915
rect 3140 -4979 3274 -4967
rect 3140 -5031 3181 -4979
rect 3233 -5031 3274 -4979
rect 3140 -5050 3274 -5031
rect 3648 -4935 3782 -4916
rect 3648 -4987 3689 -4935
rect 3741 -4987 3782 -4935
rect 3648 -4999 3782 -4987
rect 3648 -5051 3689 -4999
rect 3741 -5051 3782 -4999
rect 3648 -5070 3782 -5051
rect 388 -5134 2520 -5132
rect 388 -5168 3692 -5134
rect 388 -5170 832 -5168
rect 1012 -5192 3692 -5168
rect 4114 -5173 4153 -4673
rect 4333 -5173 4372 -4673
rect 4114 -5186 4372 -5173
rect 1012 -5200 1064 -5192
rect 442 -5224 796 -5200
rect 2420 -5210 2520 -5192
rect 4118 -5198 4368 -5186
rect 442 -5233 465 -5224
rect 442 -5260 458 -5233
rect 192 -5266 458 -5260
rect -1394 -5267 458 -5266
rect -1394 -5276 465 -5267
rect 517 -5276 529 -5224
rect 581 -5276 593 -5224
rect 645 -5276 657 -5224
rect 709 -5276 721 -5224
rect 773 -5233 796 -5224
rect 780 -5250 796 -5233
rect 1556 -5250 1818 -5226
rect 780 -5255 1818 -5250
rect 780 -5267 1597 -5255
rect 773 -5276 1597 -5267
rect -1394 -5307 1597 -5276
rect 1649 -5307 1661 -5255
rect 1713 -5307 1725 -5255
rect 1777 -5260 1818 -5255
rect 2996 -5253 3304 -5232
rect 2996 -5260 3028 -5253
rect 1777 -5262 3028 -5260
rect 1777 -5296 3025 -5262
rect 1777 -5305 3028 -5296
rect 3080 -5305 3092 -5253
rect 3144 -5305 3156 -5253
rect 3208 -5305 3220 -5253
rect 3272 -5260 3304 -5253
rect 4100 -5259 4300 -5240
rect 4100 -5260 4147 -5259
rect 3272 -5262 4147 -5260
rect 3275 -5296 4147 -5262
rect 3272 -5305 4147 -5296
rect 1777 -5307 4147 -5305
rect -1394 -5365 4147 -5307
rect 4253 -5260 4300 -5259
rect 4253 -5365 4936 -5260
rect -1394 -5654 4936 -5365
rect -1394 -5660 3350 -5654
<< via1 >>
rect 2872 631 2924 640
rect 2872 597 2873 631
rect 2873 597 2907 631
rect 2907 597 2924 631
rect 2872 588 2924 597
rect 2936 631 2988 640
rect 2936 597 2945 631
rect 2945 597 2979 631
rect 2979 597 2988 631
rect 2936 588 2988 597
rect 3000 631 3052 640
rect 3000 597 3017 631
rect 3017 597 3051 631
rect 3051 597 3052 631
rect 3000 588 3052 597
rect 3646 623 3698 632
rect 3646 589 3647 623
rect 3647 589 3681 623
rect 3681 589 3698 623
rect 3646 580 3698 589
rect 3710 623 3762 632
rect 3710 589 3719 623
rect 3719 589 3753 623
rect 3753 589 3762 623
rect 3710 580 3762 589
rect 3774 623 3826 632
rect 3774 589 3791 623
rect 3791 589 3825 623
rect 3825 589 3826 623
rect 3774 580 3826 589
rect 4412 629 4464 638
rect 4412 595 4413 629
rect 4413 595 4447 629
rect 4447 595 4464 629
rect 4412 586 4464 595
rect 4476 629 4528 638
rect 4476 595 4485 629
rect 4485 595 4519 629
rect 4519 595 4528 629
rect 4476 586 4528 595
rect 4540 629 4592 638
rect 4540 595 4557 629
rect 4557 595 4591 629
rect 4591 595 4592 629
rect 4540 586 4592 595
rect 2690 147 2742 199
rect 2690 83 2742 135
rect 2932 149 2984 201
rect 2932 85 2984 137
rect 3168 143 3220 195
rect 3168 79 3220 131
rect -1234 -1842 -1182 -1790
rect -1234 -1906 -1182 -1854
rect -1234 -1970 -1182 -1918
rect -1234 -2034 -1182 -1982
rect 1356 -953 1408 -901
rect 1356 -1017 1408 -965
rect 1356 -1081 1408 -1029
rect 1356 -1145 1408 -1093
rect 2826 -955 2878 -903
rect 2826 -1019 2878 -967
rect 2826 -1083 2878 -1031
rect 2826 -1147 2878 -1095
rect 3060 -955 3112 -903
rect 3060 -1019 3112 -967
rect 3060 -1083 3112 -1031
rect 3060 -1147 3112 -1095
rect 2254 -1760 2306 -1708
rect 2254 -1824 2306 -1772
rect 2254 -1888 2306 -1836
rect 2254 -1952 2306 -1900
rect 1916 -2280 1968 -2228
rect 1916 -2344 1968 -2292
rect 1916 -2408 1968 -2356
rect -1306 -2829 -1190 -2649
rect 884 -2855 1000 -2675
rect 1228 -3416 1280 -3364
rect 1228 -3480 1280 -3428
rect 1462 -3424 1514 -3372
rect 1462 -3488 1514 -3436
rect 1794 -3417 1846 -3365
rect 1794 -3481 1846 -3429
rect 2036 -3419 2088 -3367
rect 2036 -3483 2088 -3431
rect 3496 139 3548 191
rect 3496 75 3548 127
rect 3736 129 3788 181
rect 3736 65 3788 117
rect 3974 123 4026 175
rect 3974 59 4026 111
rect 4296 123 4348 175
rect 4296 59 4348 111
rect 4503 129 4555 181
rect 4503 65 4555 117
rect 4699 133 4751 185
rect 4699 69 4751 121
rect 3620 -2278 3672 -2226
rect 3620 -2342 3672 -2290
rect 3620 -2406 3672 -2354
rect 3854 -2284 3906 -2232
rect 3854 -2348 3906 -2296
rect 3854 -2412 3906 -2360
rect 4144 -2279 4196 -2227
rect 4144 -2343 4196 -2291
rect 4144 -2407 4196 -2355
rect 1473 -3818 1525 -3766
rect 1537 -3818 1589 -3766
rect 1601 -3818 1653 -3766
rect 1665 -3818 1717 -3766
rect 1729 -3818 1781 -3766
rect 2922 -3256 2974 -3204
rect 2922 -3320 2974 -3268
rect 3438 -3268 3490 -3216
rect 3438 -3332 3490 -3280
rect 4405 -3255 4457 -3203
rect 4405 -3319 4457 -3267
rect 4601 -3253 4653 -3201
rect 4601 -3317 4653 -3265
rect 1456 -4213 1508 -4161
rect 1456 -4277 1508 -4225
rect 1974 -4213 2026 -4161
rect 1974 -4277 2026 -4225
rect 316 -4955 368 -4903
rect 316 -5019 368 -4967
rect 316 -5083 368 -5031
rect 848 -4979 900 -4927
rect 848 -5043 900 -4991
rect 1206 -4999 1258 -4947
rect 1206 -5063 1258 -5011
rect 1716 -5009 1768 -4957
rect 1716 -5073 1768 -5021
rect 2228 -5013 2280 -4961
rect 2228 -5077 2280 -5025
rect 13087 -3602 14675 -2718
rect 2663 -4965 2715 -4913
rect 2663 -5029 2715 -4977
rect 3181 -4967 3233 -4915
rect 3181 -5031 3233 -4979
rect 3689 -4987 3741 -4935
rect 3689 -5051 3741 -4999
rect 4153 -4690 4333 -4673
rect 4153 -5156 4154 -4690
rect 4154 -5156 4332 -4690
rect 4332 -5156 4333 -4690
rect 4153 -5173 4333 -5156
rect 465 -5233 517 -5224
rect 465 -5267 492 -5233
rect 492 -5267 517 -5233
rect 465 -5276 517 -5267
rect 529 -5233 581 -5224
rect 529 -5267 530 -5233
rect 530 -5267 564 -5233
rect 564 -5267 581 -5233
rect 529 -5276 581 -5267
rect 593 -5233 645 -5224
rect 593 -5267 602 -5233
rect 602 -5267 636 -5233
rect 636 -5267 645 -5233
rect 593 -5276 645 -5267
rect 657 -5233 709 -5224
rect 657 -5267 674 -5233
rect 674 -5267 708 -5233
rect 708 -5267 709 -5233
rect 657 -5276 709 -5267
rect 721 -5233 773 -5224
rect 721 -5267 746 -5233
rect 746 -5267 773 -5233
rect 1597 -5264 1649 -5255
rect 721 -5276 773 -5267
rect 1597 -5298 1598 -5264
rect 1598 -5298 1632 -5264
rect 1632 -5298 1649 -5264
rect 1597 -5307 1649 -5298
rect 1661 -5264 1713 -5255
rect 1661 -5298 1670 -5264
rect 1670 -5298 1704 -5264
rect 1704 -5298 1713 -5264
rect 1661 -5307 1713 -5298
rect 1725 -5264 1777 -5255
rect 3028 -5262 3080 -5253
rect 1725 -5298 1742 -5264
rect 1742 -5298 1776 -5264
rect 1776 -5298 1777 -5264
rect 3028 -5296 3059 -5262
rect 3059 -5296 3080 -5262
rect 1725 -5307 1777 -5298
rect 3028 -5305 3080 -5296
rect 3092 -5262 3144 -5253
rect 3092 -5296 3097 -5262
rect 3097 -5296 3131 -5262
rect 3131 -5296 3144 -5262
rect 3092 -5305 3144 -5296
rect 3156 -5262 3208 -5253
rect 3156 -5296 3169 -5262
rect 3169 -5296 3203 -5262
rect 3203 -5296 3208 -5262
rect 3156 -5305 3208 -5296
rect 3220 -5262 3272 -5253
rect 3220 -5296 3241 -5262
rect 3241 -5296 3272 -5262
rect 3220 -5305 3272 -5296
<< metal2 >>
rect 2868 640 3056 666
rect 2868 588 2872 640
rect 2924 588 2936 640
rect 2988 588 3000 640
rect 3052 588 3056 640
rect 2868 562 3056 588
rect 3642 632 3830 658
rect 3642 580 3646 632
rect 3698 580 3710 632
rect 3762 580 3774 632
rect 3826 580 3830 632
rect 2672 199 2760 224
rect 2672 147 2690 199
rect 2742 184 2760 199
rect 2900 201 3026 562
rect 3642 554 3830 580
rect 4408 638 4596 664
rect 4408 586 4412 638
rect 4464 586 4476 638
rect 4528 586 4540 638
rect 4592 586 4596 638
rect 4408 560 4596 586
rect 2900 184 2932 201
rect 2742 149 2932 184
rect 2984 184 3026 201
rect 3150 195 3238 220
rect 3150 184 3168 195
rect 2984 149 3168 184
rect 2742 147 3168 149
rect 2672 143 3168 147
rect 3220 184 3238 195
rect 3478 191 3566 216
rect 3478 184 3496 191
rect 3220 143 3496 184
rect 2672 139 3496 143
rect 3548 184 3566 191
rect 3678 206 3804 554
rect 3678 184 3806 206
rect 3956 184 4044 200
rect 4278 184 4366 200
rect 4444 184 4570 560
rect 4688 185 4762 208
rect 4688 184 4699 185
rect 3548 181 4699 184
rect 3548 139 3736 181
rect 2672 137 3736 139
rect 2672 135 2932 137
rect 2672 83 2690 135
rect 2742 85 2932 135
rect 2984 131 3736 137
rect 2984 85 3168 131
rect 2742 83 3168 85
rect 2672 79 3168 83
rect 3220 129 3736 131
rect 3788 175 4503 181
rect 3788 129 3974 175
rect 3220 127 3974 129
rect 3220 79 3496 127
rect 2672 75 3496 79
rect 3548 123 3974 127
rect 4026 123 4296 175
rect 4348 129 4503 175
rect 4555 133 4699 181
rect 4751 133 4762 185
rect 4555 129 4762 133
rect 4348 123 4762 129
rect 3548 121 4762 123
rect 3548 117 4699 121
rect 3548 75 3736 117
rect 2672 65 3736 75
rect 3788 111 4503 117
rect 3788 65 3974 111
rect 2672 64 3974 65
rect 2672 58 2760 64
rect 2914 60 3002 64
rect 3150 54 3238 64
rect 3478 50 3566 64
rect 3718 40 3806 64
rect 3956 59 3974 64
rect 4026 64 4296 111
rect 4026 59 4044 64
rect 3956 34 4044 59
rect 4278 59 4296 64
rect 4348 65 4503 111
rect 4555 69 4699 117
rect 4751 69 4762 121
rect 4555 65 4762 69
rect 4348 64 4762 65
rect 4348 59 4366 64
rect 4278 34 4366 59
rect 4492 42 4566 64
rect 4688 46 4762 64
rect 1340 -901 1424 -866
rect 1340 -953 1356 -901
rect 1408 -950 1424 -901
rect 2810 -903 2894 -868
rect 2810 -950 2826 -903
rect 1408 -953 2826 -950
rect 1340 -955 2826 -953
rect 2878 -950 2894 -903
rect 3044 -903 3128 -868
rect 3044 -950 3060 -903
rect 2878 -955 3060 -950
rect 3112 -955 3128 -903
rect 1340 -965 3128 -955
rect 1340 -1017 1356 -965
rect 1408 -967 3128 -965
rect 1408 -1017 2826 -967
rect 1340 -1019 2826 -1017
rect 2878 -1019 3060 -967
rect 3112 -1019 3128 -967
rect 1340 -1029 3128 -1019
rect 1340 -1081 1356 -1029
rect 1408 -1031 3128 -1029
rect 1408 -1081 2826 -1031
rect 1340 -1083 2826 -1081
rect 2878 -1083 3060 -1031
rect 3112 -1083 3128 -1031
rect 1340 -1093 3128 -1083
rect 1340 -1145 1356 -1093
rect 1408 -1095 3128 -1093
rect 1408 -1104 2826 -1095
rect 1408 -1145 1424 -1104
rect 1340 -1180 1424 -1145
rect 2810 -1147 2826 -1104
rect 2878 -1104 3060 -1095
rect 2878 -1147 2894 -1104
rect 2810 -1182 2894 -1147
rect 3044 -1147 3060 -1104
rect 3112 -1147 3128 -1095
rect 3044 -1182 3128 -1147
rect 2230 -1708 2330 -1684
rect 2230 -1760 2254 -1708
rect 2306 -1760 2330 -1708
rect -1258 -1790 -1158 -1764
rect -1258 -1842 -1234 -1790
rect -1182 -1800 -1158 -1790
rect 2230 -1772 2330 -1760
rect 2230 -1800 2254 -1772
rect -1182 -1824 2254 -1800
rect 2306 -1824 2330 -1772
rect -1182 -1836 2330 -1824
rect -1182 -1842 2254 -1836
rect -1258 -1854 2254 -1842
rect -1258 -1906 -1234 -1854
rect -1182 -1888 2254 -1854
rect 2306 -1888 2330 -1836
rect -1182 -1900 2330 -1888
rect -1182 -1906 2254 -1900
rect -1258 -1918 2254 -1906
rect -1258 -1970 -1234 -1918
rect -1182 -1936 2254 -1918
rect -1182 -1970 -1158 -1936
rect -1258 -1982 -1158 -1970
rect 2230 -1952 2254 -1936
rect 2306 -1952 2330 -1900
rect 2230 -1976 2330 -1952
rect -1258 -2034 -1234 -1982
rect -1182 -2034 -1158 -1982
rect -1258 -2060 -1158 -2034
rect 1902 -2228 1982 -2188
rect 1902 -2280 1916 -2228
rect 1968 -2264 1982 -2228
rect 3606 -2226 3686 -2186
rect 3606 -2264 3620 -2226
rect 1968 -2278 3620 -2264
rect 3672 -2264 3686 -2226
rect 3840 -2232 3920 -2192
rect 3840 -2264 3854 -2232
rect 3672 -2278 3854 -2264
rect 1968 -2280 3854 -2278
rect 1902 -2284 3854 -2280
rect 3906 -2264 3920 -2232
rect 4130 -2227 4210 -2188
rect 4130 -2264 4144 -2227
rect 3906 -2279 4144 -2264
rect 4196 -2279 4210 -2227
rect 3906 -2284 4210 -2279
rect 1902 -2290 4210 -2284
rect 1902 -2292 3620 -2290
rect 1902 -2344 1916 -2292
rect 1968 -2342 3620 -2292
rect 3672 -2291 4210 -2290
rect 3672 -2296 4144 -2291
rect 3672 -2342 3854 -2296
rect 1968 -2344 3854 -2342
rect 1902 -2348 3854 -2344
rect 3906 -2343 4144 -2296
rect 4196 -2343 4210 -2291
rect 3906 -2348 4210 -2343
rect 1902 -2354 4210 -2348
rect 1902 -2356 3620 -2354
rect 1902 -2408 1916 -2356
rect 1968 -2390 3620 -2356
rect 1968 -2408 1982 -2390
rect 1902 -2448 1982 -2408
rect 3606 -2406 3620 -2390
rect 3672 -2355 4210 -2354
rect 3672 -2360 4144 -2355
rect 3672 -2390 3854 -2360
rect 3672 -2406 3686 -2390
rect 3606 -2446 3686 -2406
rect 3840 -2412 3854 -2390
rect 3906 -2390 4144 -2360
rect 3906 -2412 3920 -2390
rect 3840 -2452 3920 -2412
rect 4130 -2407 4144 -2390
rect 4196 -2407 4210 -2355
rect 4130 -2446 4210 -2407
rect -1308 -2649 -1188 -2610
rect -1308 -2829 -1306 -2649
rect -1190 -2668 -1188 -2649
rect 882 -2668 1002 -2636
rect -1190 -2675 1002 -2668
rect -1190 -2829 884 -2675
rect -1308 -2848 884 -2829
rect -1308 -2868 -1188 -2848
rect 882 -2855 884 -2848
rect 1000 -2855 1002 -2675
rect 882 -2894 1002 -2855
rect 13058 -2692 14704 -2682
rect 13058 -2718 13093 -2692
rect 14669 -2718 14704 -2692
rect 13058 -3018 13087 -2718
rect 11890 -3048 13087 -3018
rect 2870 -3050 4152 -3048
rect 4314 -3050 13087 -3048
rect 2870 -3201 13087 -3050
rect 2870 -3203 4601 -3201
rect 2870 -3204 4405 -3203
rect 2870 -3256 2922 -3204
rect 2974 -3216 4405 -3204
rect 2974 -3256 3438 -3216
rect 2870 -3268 3438 -3256
rect 3490 -3255 4405 -3216
rect 4457 -3253 4601 -3203
rect 4653 -3253 13087 -3201
rect 4457 -3255 13087 -3253
rect 3490 -3265 13087 -3255
rect 3490 -3267 4601 -3265
rect 3490 -3268 4405 -3267
rect 2870 -3320 2922 -3268
rect 2974 -3280 4405 -3268
rect 2974 -3320 3438 -3280
rect 1210 -3364 1298 -3326
rect 1210 -3416 1228 -3364
rect 1280 -3384 1298 -3364
rect 1444 -3372 1532 -3334
rect 1444 -3384 1462 -3372
rect 1280 -3416 1462 -3384
rect 1210 -3424 1462 -3416
rect 1514 -3384 1532 -3372
rect 1784 -3365 1856 -3330
rect 2870 -3332 3438 -3320
rect 3490 -3319 4405 -3280
rect 4457 -3317 4601 -3267
rect 4653 -3317 13087 -3265
rect 4457 -3319 13087 -3317
rect 3490 -3332 13087 -3319
rect 1784 -3384 1794 -3365
rect 1514 -3417 1794 -3384
rect 1846 -3384 1856 -3365
rect 2026 -3367 2098 -3332
rect 2026 -3384 2036 -3367
rect 1846 -3417 2036 -3384
rect 1514 -3419 2036 -3417
rect 2088 -3419 2098 -3367
rect 2870 -3382 13087 -3332
rect 2870 -3388 12342 -3382
rect 2870 -3396 4152 -3388
rect 4314 -3396 12342 -3388
rect 1514 -3424 2098 -3419
rect 1210 -3428 2098 -3424
rect 1210 -3480 1228 -3428
rect 1280 -3429 2098 -3428
rect 1280 -3436 1794 -3429
rect 1280 -3480 1462 -3436
rect 1210 -3488 1462 -3480
rect 1514 -3481 1794 -3436
rect 1846 -3431 2098 -3429
rect 1846 -3481 2036 -3431
rect 1514 -3483 2036 -3481
rect 2088 -3483 2098 -3431
rect 1514 -3488 2098 -3483
rect 1210 -3490 2098 -3488
rect 1210 -3518 1298 -3490
rect 1444 -3526 1532 -3490
rect 1784 -3516 1856 -3490
rect 1906 -3518 2098 -3490
rect 1452 -3736 1802 -3726
rect 1132 -3766 1802 -3736
rect 1132 -3818 1473 -3766
rect 1525 -3818 1537 -3766
rect 1589 -3818 1601 -3766
rect 1653 -3818 1665 -3766
rect 1717 -3818 1729 -3766
rect 1781 -3818 1802 -3766
rect 1132 -3848 1802 -3818
rect 296 -4903 388 -4892
rect 296 -4955 316 -4903
rect 368 -4906 388 -4903
rect 368 -4927 930 -4906
rect 368 -4955 848 -4927
rect 296 -4967 848 -4955
rect 296 -5019 316 -4967
rect 368 -4979 848 -4967
rect 900 -4934 930 -4927
rect 1132 -4934 1290 -3848
rect 1452 -3858 1802 -3848
rect 1430 -4161 1534 -4134
rect 1430 -4213 1456 -4161
rect 1508 -4164 1534 -4161
rect 1906 -4161 2070 -3518
rect 13058 -3602 13087 -3382
rect 14675 -3602 14704 -2718
rect 13058 -3628 13093 -3602
rect 14669 -3628 14704 -3602
rect 13058 -3638 14704 -3628
rect 1906 -4164 1974 -4161
rect 1508 -4213 1974 -4164
rect 2026 -4174 2070 -4161
rect 2026 -4213 2052 -4174
rect 1430 -4225 2052 -4213
rect 1430 -4277 1456 -4225
rect 1508 -4277 1974 -4225
rect 2026 -4277 2052 -4225
rect 1430 -4278 2052 -4277
rect 1430 -4304 1534 -4278
rect 1948 -4304 2052 -4278
rect 4124 -4673 4362 -4650
rect 4124 -4695 4153 -4673
rect 4333 -4695 4362 -4673
rect 2632 -4913 2746 -4884
rect 2632 -4918 2663 -4913
rect 900 -4947 1290 -4934
rect 900 -4979 1206 -4947
rect 368 -4991 1206 -4979
rect 368 -5019 848 -4991
rect 296 -5031 848 -5019
rect 296 -5083 316 -5031
rect 368 -5043 848 -5031
rect 900 -4999 1206 -4991
rect 1258 -4960 1290 -4947
rect 1690 -4957 1794 -4930
rect 1690 -4960 1716 -4957
rect 1258 -4999 1716 -4960
rect 900 -5009 1716 -4999
rect 1768 -4960 1794 -4957
rect 2120 -4960 2663 -4918
rect 1768 -4961 2663 -4960
rect 1768 -5009 2228 -4961
rect 900 -5011 2228 -5009
rect 900 -5043 1206 -5011
rect 368 -5054 1206 -5043
rect 368 -5068 930 -5054
rect 1180 -5063 1206 -5054
rect 1258 -5013 2228 -5011
rect 2280 -4965 2663 -4961
rect 2715 -4918 2746 -4913
rect 3150 -4915 3264 -4886
rect 2715 -4924 2788 -4918
rect 3150 -4924 3181 -4915
rect 2715 -4965 3181 -4924
rect 2280 -4967 3181 -4965
rect 3233 -4924 3264 -4915
rect 3658 -4924 3772 -4906
rect 3233 -4935 3772 -4924
rect 3233 -4967 3689 -4935
rect 2280 -4977 3689 -4967
rect 2280 -5013 2663 -4977
rect 1258 -5021 2663 -5013
rect 1258 -5063 1716 -5021
rect 368 -5083 388 -5068
rect 296 -5094 388 -5083
rect 554 -5196 666 -5068
rect 1180 -5073 1716 -5063
rect 1768 -5025 2663 -5021
rect 1768 -5073 2228 -5025
rect 1180 -5077 2228 -5073
rect 2280 -5029 2663 -5025
rect 2715 -4979 3689 -4977
rect 2715 -5029 3181 -4979
rect 2280 -5031 3181 -5029
rect 3233 -4987 3689 -4979
rect 3741 -4987 3772 -4935
rect 3233 -4999 3772 -4987
rect 3233 -5031 3689 -4999
rect 2280 -5040 3689 -5031
rect 2280 -5076 2788 -5040
rect 2280 -5077 2306 -5076
rect 1180 -5082 2306 -5077
rect 1180 -5090 1284 -5082
rect 1610 -5100 1794 -5082
rect 454 -5224 784 -5196
rect 1610 -5222 1778 -5100
rect 2202 -5104 2306 -5082
rect 454 -5276 465 -5224
rect 517 -5276 529 -5224
rect 581 -5276 593 -5224
rect 645 -5276 657 -5224
rect 709 -5276 721 -5224
rect 773 -5276 784 -5224
rect 454 -5304 784 -5276
rect 1568 -5255 1806 -5222
rect 3130 -5228 3278 -5040
rect 3658 -5051 3689 -5040
rect 3741 -5051 3772 -4999
rect 3658 -5080 3772 -5051
rect 4124 -5151 4135 -4695
rect 4351 -5151 4362 -4695
rect 4124 -5173 4153 -5151
rect 4333 -5173 4362 -5151
rect 4124 -5196 4362 -5173
rect 1568 -5307 1597 -5255
rect 1649 -5307 1661 -5255
rect 1713 -5307 1725 -5255
rect 1777 -5307 1806 -5255
rect 1568 -5340 1806 -5307
rect 3008 -5253 3292 -5228
rect 3008 -5305 3028 -5253
rect 3080 -5305 3092 -5253
rect 3144 -5305 3156 -5253
rect 3208 -5305 3220 -5253
rect 3272 -5305 3292 -5253
rect 3008 -5330 3292 -5305
<< via2 >>
rect 13093 -2718 14669 -2692
rect 13093 -3602 14669 -2718
rect 13093 -3628 14669 -3602
rect 4135 -5151 4153 -4695
rect 4153 -5151 4333 -4695
rect 4333 -5151 4351 -4695
<< metal3 >>
rect 13048 -2692 14714 -2687
rect 13048 -2728 13093 -2692
rect 14669 -2728 14714 -2692
rect 13048 -3592 13089 -2728
rect 14673 -3592 14714 -2728
rect 13048 -3628 13093 -3592
rect 14669 -3628 14714 -3592
rect 13048 -3633 14714 -3628
rect 4114 -4691 4372 -4655
rect 4114 -5155 4131 -4691
rect 4355 -5155 4372 -4691
rect 4114 -5191 4372 -5155
<< via3 >>
rect 13089 -3592 13093 -2728
rect 13093 -3592 14669 -2728
rect 14669 -3592 14673 -2728
rect 4131 -4695 4355 -4691
rect 4131 -5151 4135 -4695
rect 4135 -5151 4351 -4695
rect 4351 -5151 4355 -4695
rect 4131 -5155 4355 -5151
<< metal4 >>
rect 11412 -2691 13096 -2690
rect 11412 -2728 14705 -2691
rect 11412 -3592 13089 -2728
rect 14673 -3592 14705 -2728
rect 11412 -3628 14705 -3592
rect 13057 -3629 14705 -3628
rect 3894 -4691 5174 -4528
rect 3894 -5155 4131 -4691
rect 4355 -5155 5174 -4691
rect 3894 -5214 5174 -5155
use sky130_fd_pr__cap_mim_m3_1_ALHCBP  sky130_fd_pr__cap_mim_m3_1_ALHCBP_0
timestamp 1725256412
transform 1 0 8278 0 1 -2308
box -3186 -3040 3186 3040
use sky130_fd_pr__nfet_01v8_24RZ45  XM9
timestamp 1725256412
transform 1 0 3203 0 1 -4106
box -673 -1200 673 1200
use sky130_fd_pr__pfet_01v8_R7N38B  XM10
timestamp 1725256412
transform 1 0 4529 0 1 -1475
box -363 -2119 363 2119
use sky130_fd_pr__pfet_01v8_Q9ENJR  XM11
timestamp 1725256412
transform 1 0 2957 0 1 -1075
box -403 -1719 403 1719
use sky130_fd_pr__nfet_01v8_7PL8E9  XM12
timestamp 1725256412
transform 1 0 1941 0 1 -2100
box -275 -1700 275 1700
use sky130_fd_pr__nfet_01v8_7PL8E9  XM13
timestamp 1725256412
transform 1 0 1371 0 1 -2100
box -275 -1700 275 1700
use sky130_fd_pr__nfet_01v8_4G38HM  XM14
timestamp 1725256412
transform 1 0 1741 0 1 -4596
box -673 -700 673 700
use sky130_fd_pr__pfet_01v8_Q9ENJR  XM15
timestamp 1725256412
transform 1 0 3763 0 1 -1075
box -403 -1719 403 1719
use sky130_fd_pr__nfet_01v8_JCA7Y6  XM16
timestamp 1725256412
transform 1 0 617 0 1 -4982
box -415 -300 415 300
use sky130_fd_pr__res_high_po_0p69_UD9NEZ  XR1
timestamp 1725256412
transform 1 0 4231 0 1 -4544
box -225 -762 225 762
use sky130_fd_pr__res_high_po_0p35_BQ2QQJ  XR2
timestamp 1725256412
transform 1 0 407 0 1 -2192
box -191 -2472 191 2472
use sky130_fd_pr__res_high_po_0p35_BQ2QQJ  XR3
timestamp 1725256412
transform 1 0 7 0 1 -2192
box -191 -2472 191 2472
use sky130_fd_pr__res_high_po_0p35_BQ2QQJ  XR4
timestamp 1725256412
transform 1 0 -395 0 1 -2192
box -191 -2472 191 2472
use sky130_fd_pr__res_high_po_0p35_BQ2QQJ  XR5
timestamp 1725256412
transform 1 0 -795 0 1 -2192
box -191 -2472 191 2472
use sky130_fd_pr__res_high_po_0p35_BQ2QQJ  XR14
timestamp 1725256412
transform 1 0 809 0 1 -2192
box -191 -2472 191 2472
<< labels >>
flabel metal1 s 3632 658 3832 858 0 FreeSans 400 0 0 0 VDD
port 1 nsew
flabel metal1 s -1404 -2812 -1204 -2612 0 FreeSans 400 0 0 0 INP
port 2 nsew
flabel metal1 s -1306 -2000 -1106 -1800 0 FreeSans 400 0 0 0 INN
port 3 nsew
flabel metal2 s 13622 -3274 13822 -3074 0 FreeSans 400 0 0 0 VOUT
port 4 nsew
flabel metal1 s 1052 -5628 1252 -5428 0 FreeSans 400 0 0 0 VSS
port 5 nsew
<< end >>
