magic
tech sky130A
magscale 1 2
timestamp 1725467580
<< nmoslvt >>
rect -3403 -431 -2603 369
rect -2545 -431 -1745 369
rect -1687 -431 -887 369
rect -829 -431 -29 369
rect 29 -431 829 369
rect 887 -431 1687 369
rect 1745 -431 2545 369
rect 2603 -431 3403 369
<< ndiff >>
rect -3461 357 -3403 369
rect -3461 -419 -3449 357
rect -3415 -419 -3403 357
rect -3461 -431 -3403 -419
rect -2603 357 -2545 369
rect -2603 -419 -2591 357
rect -2557 -419 -2545 357
rect -2603 -431 -2545 -419
rect -1745 357 -1687 369
rect -1745 -419 -1733 357
rect -1699 -419 -1687 357
rect -1745 -431 -1687 -419
rect -887 357 -829 369
rect -887 -419 -875 357
rect -841 -419 -829 357
rect -887 -431 -829 -419
rect -29 357 29 369
rect -29 -419 -17 357
rect 17 -419 29 357
rect -29 -431 29 -419
rect 829 357 887 369
rect 829 -419 841 357
rect 875 -419 887 357
rect 829 -431 887 -419
rect 1687 357 1745 369
rect 1687 -419 1699 357
rect 1733 -419 1745 357
rect 1687 -431 1745 -419
rect 2545 357 2603 369
rect 2545 -419 2557 357
rect 2591 -419 2603 357
rect 2545 -431 2603 -419
rect 3403 357 3461 369
rect 3403 -419 3415 357
rect 3449 -419 3461 357
rect 3403 -431 3461 -419
<< ndiffc >>
rect -3449 -419 -3415 357
rect -2591 -419 -2557 357
rect -1733 -419 -1699 357
rect -875 -419 -841 357
rect -17 -419 17 357
rect 841 -419 875 357
rect 1699 -419 1733 357
rect 2557 -419 2591 357
rect 3415 -419 3449 357
<< poly >>
rect -3403 441 -2603 457
rect -3403 407 -3387 441
rect -2619 407 -2603 441
rect -3403 369 -2603 407
rect -2545 441 -1745 457
rect -2545 407 -2529 441
rect -1761 407 -1745 441
rect -2545 369 -1745 407
rect -1687 441 -887 457
rect -1687 407 -1671 441
rect -903 407 -887 441
rect -1687 369 -887 407
rect -829 441 -29 457
rect -829 407 -813 441
rect -45 407 -29 441
rect -829 369 -29 407
rect 29 441 829 457
rect 29 407 45 441
rect 813 407 829 441
rect 29 369 829 407
rect 887 441 1687 457
rect 887 407 903 441
rect 1671 407 1687 441
rect 887 369 1687 407
rect 1745 441 2545 457
rect 1745 407 1761 441
rect 2529 407 2545 441
rect 1745 369 2545 407
rect 2603 441 3403 457
rect 2603 407 2619 441
rect 3387 407 3403 441
rect 2603 369 3403 407
rect -3403 -457 -2603 -431
rect -2545 -457 -1745 -431
rect -1687 -457 -887 -431
rect -829 -457 -29 -431
rect 29 -457 829 -431
rect 887 -457 1687 -431
rect 1745 -457 2545 -431
rect 2603 -457 3403 -431
<< polycont >>
rect -3387 407 -2619 441
rect -2529 407 -1761 441
rect -1671 407 -903 441
rect -813 407 -45 441
rect 45 407 813 441
rect 903 407 1671 441
rect 1761 407 2529 441
rect 2619 407 3387 441
<< locali >>
rect -3403 407 -3387 441
rect -2619 407 -2603 441
rect -2545 407 -2529 441
rect -1761 407 -1745 441
rect -1687 407 -1671 441
rect -903 407 -887 441
rect -829 407 -813 441
rect -45 407 -29 441
rect 29 407 45 441
rect 813 407 829 441
rect 887 407 903 441
rect 1671 407 1687 441
rect 1745 407 1761 441
rect 2529 407 2545 441
rect 2603 407 2619 441
rect 3387 407 3403 441
rect -3449 357 -3415 373
rect -3449 -435 -3415 -419
rect -2591 357 -2557 373
rect -2591 -435 -2557 -419
rect -1733 357 -1699 373
rect -1733 -435 -1699 -419
rect -875 357 -841 373
rect -875 -435 -841 -419
rect -17 357 17 373
rect -17 -435 17 -419
rect 841 357 875 373
rect 841 -435 875 -419
rect 1699 357 1733 373
rect 1699 -435 1733 -419
rect 2557 357 2591 373
rect 2557 -435 2591 -419
rect 3415 357 3449 373
rect 3415 -435 3449 -419
<< viali >>
rect -3387 407 -2619 441
rect -2529 407 -1761 441
rect -1671 407 -903 441
rect -813 407 -45 441
rect 45 407 813 441
rect 903 407 1671 441
rect 1761 407 2529 441
rect 2619 407 3387 441
rect -3449 107 -3415 340
rect -2591 -402 -2557 -169
rect -1733 107 -1699 340
rect -875 -402 -841 -169
rect -17 107 17 340
rect 841 -402 875 -169
rect 1699 107 1733 340
rect 2557 -402 2591 -169
rect 3415 107 3449 340
<< metal1 >>
rect -3399 441 -2607 447
rect -3399 407 -3387 441
rect -2619 407 -2607 441
rect -3399 401 -2607 407
rect -2541 441 -1749 447
rect -2541 407 -2529 441
rect -1761 407 -1749 441
rect -2541 401 -1749 407
rect -1683 441 -891 447
rect -1683 407 -1671 441
rect -903 407 -891 441
rect -1683 401 -891 407
rect -825 441 -33 447
rect -825 407 -813 441
rect -45 407 -33 441
rect -825 401 -33 407
rect 33 441 825 447
rect 33 407 45 441
rect 813 407 825 441
rect 33 401 825 407
rect 891 441 1683 447
rect 891 407 903 441
rect 1671 407 1683 441
rect 891 401 1683 407
rect 1749 441 2541 447
rect 1749 407 1761 441
rect 2529 407 2541 441
rect 1749 401 2541 407
rect 2607 441 3399 447
rect 2607 407 2619 441
rect 3387 407 3399 441
rect 2607 401 3399 407
rect -3455 340 -3409 352
rect -3455 107 -3449 340
rect -3415 107 -3409 340
rect -3455 95 -3409 107
rect -1739 340 -1693 352
rect -1739 107 -1733 340
rect -1699 107 -1693 340
rect -1739 95 -1693 107
rect -23 340 23 352
rect -23 107 -17 340
rect 17 107 23 340
rect -23 95 23 107
rect 1693 340 1739 352
rect 1693 107 1699 340
rect 1733 107 1739 340
rect 1693 95 1739 107
rect 3409 340 3455 352
rect 3409 107 3415 340
rect 3449 107 3455 340
rect 3409 95 3455 107
rect -2597 -169 -2551 -157
rect -2597 -402 -2591 -169
rect -2557 -402 -2551 -169
rect -2597 -414 -2551 -402
rect -881 -169 -835 -157
rect -881 -402 -875 -169
rect -841 -402 -835 -169
rect -881 -414 -835 -402
rect 835 -169 881 -157
rect 835 -402 841 -169
rect 875 -402 881 -169
rect 835 -414 881 -402
rect 2551 -169 2597 -157
rect 2551 -402 2557 -169
rect 2591 -402 2597 -169
rect 2551 -414 2597 -402
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 4 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
