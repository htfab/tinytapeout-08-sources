magic
tech sky130A
magscale 1 2
timestamp 1725467580
<< nmoslvt >>
rect -3403 -369 -2603 431
rect -2545 -369 -1745 431
rect -1687 -369 -887 431
rect -829 -369 -29 431
rect 29 -369 829 431
rect 887 -369 1687 431
rect 1745 -369 2545 431
rect 2603 -369 3403 431
<< ndiff >>
rect -3461 419 -3403 431
rect -3461 -357 -3449 419
rect -3415 -357 -3403 419
rect -3461 -369 -3403 -357
rect -2603 419 -2545 431
rect -2603 -357 -2591 419
rect -2557 -357 -2545 419
rect -2603 -369 -2545 -357
rect -1745 419 -1687 431
rect -1745 -357 -1733 419
rect -1699 -357 -1687 419
rect -1745 -369 -1687 -357
rect -887 419 -829 431
rect -887 -357 -875 419
rect -841 -357 -829 419
rect -887 -369 -829 -357
rect -29 419 29 431
rect -29 -357 -17 419
rect 17 -357 29 419
rect -29 -369 29 -357
rect 829 419 887 431
rect 829 -357 841 419
rect 875 -357 887 419
rect 829 -369 887 -357
rect 1687 419 1745 431
rect 1687 -357 1699 419
rect 1733 -357 1745 419
rect 1687 -369 1745 -357
rect 2545 419 2603 431
rect 2545 -357 2557 419
rect 2591 -357 2603 419
rect 2545 -369 2603 -357
rect 3403 419 3461 431
rect 3403 -357 3415 419
rect 3449 -357 3461 419
rect 3403 -369 3461 -357
<< ndiffc >>
rect -3449 -357 -3415 419
rect -2591 -357 -2557 419
rect -1733 -357 -1699 419
rect -875 -357 -841 419
rect -17 -357 17 419
rect 841 -357 875 419
rect 1699 -357 1733 419
rect 2557 -357 2591 419
rect 3415 -357 3449 419
<< poly >>
rect -3403 431 -2603 457
rect -2545 431 -1745 457
rect -1687 431 -887 457
rect -829 431 -29 457
rect 29 431 829 457
rect 887 431 1687 457
rect 1745 431 2545 457
rect 2603 431 3403 457
rect -3403 -407 -2603 -369
rect -3403 -441 -3387 -407
rect -2619 -441 -2603 -407
rect -3403 -457 -2603 -441
rect -2545 -407 -1745 -369
rect -2545 -441 -2529 -407
rect -1761 -441 -1745 -407
rect -2545 -457 -1745 -441
rect -1687 -407 -887 -369
rect -1687 -441 -1671 -407
rect -903 -441 -887 -407
rect -1687 -457 -887 -441
rect -829 -407 -29 -369
rect -829 -441 -813 -407
rect -45 -441 -29 -407
rect -829 -457 -29 -441
rect 29 -407 829 -369
rect 29 -441 45 -407
rect 813 -441 829 -407
rect 29 -457 829 -441
rect 887 -407 1687 -369
rect 887 -441 903 -407
rect 1671 -441 1687 -407
rect 887 -457 1687 -441
rect 1745 -407 2545 -369
rect 1745 -441 1761 -407
rect 2529 -441 2545 -407
rect 1745 -457 2545 -441
rect 2603 -407 3403 -369
rect 2603 -441 2619 -407
rect 3387 -441 3403 -407
rect 2603 -457 3403 -441
<< polycont >>
rect -3387 -441 -2619 -407
rect -2529 -441 -1761 -407
rect -1671 -441 -903 -407
rect -813 -441 -45 -407
rect 45 -441 813 -407
rect 903 -441 1671 -407
rect 1761 -441 2529 -407
rect 2619 -441 3387 -407
<< locali >>
rect -3449 419 -3415 435
rect -3449 -373 -3415 -357
rect -2591 419 -2557 435
rect -2591 -373 -2557 -357
rect -1733 419 -1699 435
rect -1733 -373 -1699 -357
rect -875 419 -841 435
rect -875 -373 -841 -357
rect -17 419 17 435
rect -17 -373 17 -357
rect 841 419 875 435
rect 841 -373 875 -357
rect 1699 419 1733 435
rect 1699 -373 1733 -357
rect 2557 419 2591 435
rect 2557 -373 2591 -357
rect 3415 419 3449 435
rect 3415 -373 3449 -357
rect -3403 -441 -3387 -407
rect -2619 -441 -2603 -407
rect -2545 -441 -2529 -407
rect -1761 -441 -1745 -407
rect -1687 -441 -1671 -407
rect -903 -441 -887 -407
rect -829 -441 -813 -407
rect -45 -441 -29 -407
rect 29 -441 45 -407
rect 813 -441 829 -407
rect 887 -441 903 -407
rect 1671 -441 1687 -407
rect 1745 -441 1761 -407
rect 2529 -441 2545 -407
rect 2603 -441 2619 -407
rect 3387 -441 3403 -407
<< viali >>
rect -3449 169 -3415 402
rect -2591 -340 -2557 -107
rect -1733 169 -1699 402
rect -875 -340 -841 -107
rect -17 169 17 402
rect 841 -340 875 -107
rect 1699 169 1733 402
rect 2557 -340 2591 -107
rect 3415 169 3449 402
rect -3387 -441 -2619 -407
rect -2529 -441 -1761 -407
rect -1671 -441 -903 -407
rect -813 -441 -45 -407
rect 45 -441 813 -407
rect 903 -441 1671 -407
rect 1761 -441 2529 -407
rect 2619 -441 3387 -407
<< metal1 >>
rect -3455 402 -3409 414
rect -3455 169 -3449 402
rect -3415 169 -3409 402
rect -3455 157 -3409 169
rect -1739 402 -1693 414
rect -1739 169 -1733 402
rect -1699 169 -1693 402
rect -1739 157 -1693 169
rect -23 402 23 414
rect -23 169 -17 402
rect 17 169 23 402
rect -23 157 23 169
rect 1693 402 1739 414
rect 1693 169 1699 402
rect 1733 169 1739 402
rect 1693 157 1739 169
rect 3409 402 3455 414
rect 3409 169 3415 402
rect 3449 169 3455 402
rect 3409 157 3455 169
rect -2597 -107 -2551 -95
rect -2597 -340 -2591 -107
rect -2557 -340 -2551 -107
rect -2597 -352 -2551 -340
rect -881 -107 -835 -95
rect -881 -340 -875 -107
rect -841 -340 -835 -107
rect -881 -352 -835 -340
rect 835 -107 881 -95
rect 835 -340 841 -107
rect 875 -340 881 -107
rect 835 -352 881 -340
rect 2551 -107 2597 -95
rect 2551 -340 2557 -107
rect 2591 -340 2597 -107
rect 2551 -352 2597 -340
rect -3399 -407 -2607 -401
rect -3399 -441 -3387 -407
rect -2619 -441 -2607 -407
rect -3399 -447 -2607 -441
rect -2541 -407 -1749 -401
rect -2541 -441 -2529 -407
rect -1761 -441 -1749 -407
rect -2541 -447 -1749 -441
rect -1683 -407 -891 -401
rect -1683 -441 -1671 -407
rect -903 -441 -891 -407
rect -1683 -447 -891 -441
rect -825 -407 -33 -401
rect -825 -441 -813 -407
rect -45 -441 -33 -407
rect -825 -447 -33 -441
rect 33 -407 825 -401
rect 33 -441 45 -407
rect 813 -441 825 -407
rect 33 -447 825 -441
rect 891 -407 1683 -401
rect 891 -441 903 -407
rect 1671 -441 1683 -407
rect 891 -447 1683 -441
rect 1749 -407 2541 -401
rect 1749 -441 1761 -407
rect 2529 -441 2541 -407
rect 1749 -447 2541 -441
rect 2607 -407 3399 -401
rect 2607 -441 2619 -407
rect 3387 -441 3399 -407
rect 2607 -447 3399 -441
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 4 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc +30 viadrn -30 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
