magic
tech sky130A
magscale 1 2
timestamp 1725442979
<< locali >>
rect 630 390 1370 450
rect 630 310 830 390
rect 1170 310 1370 390
rect 630 280 1370 310
rect 630 -210 830 280
rect 1170 -210 1370 280
rect 630 -780 840 -300
rect 1160 -780 1370 -300
rect 630 -810 1370 -780
rect 630 -890 830 -810
rect 1170 -890 1370 -810
rect 630 -950 1370 -890
<< viali >>
rect 830 310 1170 390
rect 830 -890 1170 -810
<< metal1 >>
rect 630 400 830 450
rect 1170 400 1370 450
rect 630 390 1370 400
rect 630 310 830 390
rect 1170 310 1370 390
rect 630 300 1370 310
rect 630 250 830 300
rect 930 -30 980 300
rect 1170 250 1370 300
rect 1030 10 1070 170
rect 1030 -30 1180 10
rect 630 -230 830 -160
rect 970 -230 1030 -70
rect 630 -280 1030 -230
rect 630 -360 830 -280
rect 970 -440 1030 -280
rect 1140 -160 1180 -30
rect 1140 -360 1370 -160
rect 1140 -470 1180 -360
rect 630 -800 830 -750
rect 930 -800 980 -470
rect 1020 -510 1180 -470
rect 1020 -670 1070 -510
rect 1170 -800 1370 -750
rect 630 -810 1370 -800
rect 630 -890 830 -810
rect 1170 -890 1370 -810
rect 630 -900 1370 -890
rect 630 -950 830 -900
rect 1170 -950 1370 -900
use sky130_fd_pr__nfet_01v8_64Z3AY  XM1
timestamp 1725442979
transform 1 0 1001 0 1 -541
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_LGS3BL  XM2
timestamp 1725442979
transform 1 0 1001 0 1 34
box -211 -284 211 284
<< labels >>
flabel metal1 630 250 830 450 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 630 -360 830 -160 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 1170 -360 1370 -160 0 FreeSans 256 0 0 0 Vout
port 2 nsew
flabel metal1 630 -950 830 -750 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
